
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCRSL, SGE, 
   SLE, SNE, aluNOP);
attribute ENUM_ENCODING of aluOp : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010 1011";

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_add_1_DW01_add_3 is

   port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (29 downto 0);  CO : out std_logic);

end ALU_N32_DW01_add_1_DW01_add_3;

architecture SYN_cla of ALU_N32_DW01_add_1_DW01_add_3 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, SUM_25_port, 
      SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, 
      SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, n1, n2, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n398, n399, n400, 
      n401, SUM_14_port, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415 : std_logic;

begin
   SUM <= ( SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, SUM_25_port, 
      SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, 
      SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, 
      SUM_14_port, A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), 
      A(4), A(3), A(2), A(1), A(0) );
   
   U6 : XOR2_X1 port map( A => n37, B => n1, Z => SUM_27_port);
   U8 : XOR2_X1 port map( A => n41, B => n2, Z => SUM_25_port);
   U24 : XOR2_X1 port map( A => n21, B => n22, Z => SUM_29_port);
   U27 : XOR2_X1 port map( A => n23, B => n26, Z => SUM_28_port);
   U47 : XOR2_X1 port map( A => n43, B => n44, Z => SUM_24_port);
   U71 : XOR2_X1 port map( A => n63, B => n64, Z => SUM_20_port);
   U100 : XOR2_X1 port map( A => n86, B => n88, Z => SUM_15_port);
   U9 : XOR2_X1 port map( A => n80, B => n90, Z => SUM_17_port);
   U46 : XOR2_X1 port map( A => n60, B => n91, Z => SUM_21_port);
   U2 : OAI21_X1 port map( B1 => n80, B2 => n72, A => n74, ZN => n77);
   U3 : NAND2_X1 port map( A1 => n404, A2 => n74, ZN => n90);
   U4 : NOR2_X1 port map( A1 => n69, A2 => n403, ZN => n80);
   U5 : NOR2_X1 port map( A1 => n49, A2 => n413, ZN => n60);
   U7 : NOR2_X1 port map( A1 => n31, A2 => n409, ZN => n41);
   U10 : INV_X1 port map( A => n73, ZN => n403);
   U11 : INV_X1 port map( A => n72, ZN => n404);
   U12 : NOR2_X1 port map( A1 => B(17), A2 => A(17), ZN => n72);
   U13 : OAI21_X1 port map( B1 => n60, B2 => n52, A => n54, ZN => n57);
   U14 : OAI21_X1 port map( B1 => n41, B2 => n34, A => n36, ZN => n38);
   U15 : NOR2_X1 port map( A1 => n62, A2 => n413, ZN => n64);
   U16 : NAND2_X1 port map( A1 => n412, A2 => n54, ZN => n91);
   U17 : NOR2_X1 port map( A1 => n42, A2 => n409, ZN => n44);
   U18 : NAND2_X1 port map( A1 => n408, A2 => n36, ZN => n2);
   U19 : NAND2_X1 port map( A1 => n406, A2 => n29, ZN => n1);
   U20 : AOI21_X1 port map( B1 => n38, B2 => n32, A => n407, ZN => n37);
   U21 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => n26);
   U22 : OAI211_X1 port map( C1 => n65, C2 => n66, A => n67, B => n68, ZN => 
                           n63);
   U23 : NAND4_X1 port map( A1 => n69, A2 => n404, A3 => n70, A4 => n414, ZN =>
                           n68);
   U25 : AOI21_X1 port map( B1 => n70, B2 => n71, A => n405, ZN => n65);
   U26 : OAI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n71);
   U28 : OAI211_X1 port map( C1 => n45, C2 => n46, A => n47, B => n48, ZN => 
                           n43);
   U29 : NAND4_X1 port map( A1 => n49, A2 => n412, A3 => n50, A4 => n410, ZN =>
                           n48);
   U30 : AOI21_X1 port map( B1 => n50, B2 => n51, A => n411, ZN => n45);
   U31 : OAI21_X1 port map( B1 => n52, B2 => n53, A => n54, ZN => n51);
   U32 : OAI211_X1 port map( C1 => n27, C2 => n28, A => n29, B => n30, ZN => 
                           n23);
   U33 : NAND4_X1 port map( A1 => n31, A2 => n408, A3 => n32, A4 => n406, ZN =>
                           n30);
   U34 : AOI21_X1 port map( B1 => n32, B2 => n33, A => n407, ZN => n27);
   U35 : OAI21_X1 port map( B1 => n34, B2 => n35, A => n36, ZN => n33);
   U36 : NOR2_X1 port map( A1 => B(16), A2 => A(16), ZN => n82);
   U37 : NOR2_X1 port map( A1 => B(15), A2 => A(15), ZN => n85);
   U38 : NOR2_X1 port map( A1 => n401, A2 => n82, ZN => n69);
   U39 : NOR2_X1 port map( A1 => n400, A2 => n62, ZN => n49);
   U40 : INV_X1 port map( A => n63, ZN => n400);
   U41 : NOR2_X1 port map( A1 => n399, A2 => n42, ZN => n31);
   U42 : INV_X1 port map( A => n43, ZN => n399);
   U43 : XNOR2_X1 port map( A => n79, B => n77, ZN => SUM_18_port);
   U44 : NAND2_X1 port map( A1 => n78, A2 => n70, ZN => n79);
   U45 : XNOR2_X1 port map( A => n59, B => n57, ZN => SUM_22_port);
   U48 : NAND2_X1 port map( A1 => n58, A2 => n50, ZN => n59);
   U49 : XNOR2_X1 port map( A => n40, B => n38, ZN => SUM_26_port);
   U50 : NAND2_X1 port map( A1 => n39, A2 => n32, ZN => n40);
   U51 : XNOR2_X1 port map( A => n401, B => n83, ZN => SUM_16_port);
   U52 : NOR2_X1 port map( A1 => n82, A2 => n403, ZN => n83);
   U53 : XNOR2_X1 port map( A => n75, B => n76, ZN => SUM_19_port);
   U54 : AND2_X1 port map( A1 => n414, A2 => n67, ZN => n76);
   U55 : AOI21_X1 port map( B1 => n77, B2 => n70, A => n405, ZN => n75);
   U56 : XNOR2_X1 port map( A => n55, B => n56, ZN => SUM_23_port);
   U57 : AND2_X1 port map( A1 => n410, A2 => n47, ZN => n56);
   U58 : AOI21_X1 port map( B1 => n57, B2 => n50, A => n411, ZN => n55);
   U59 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => n74);
   U60 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n73);
   U61 : NAND2_X1 port map( A1 => B(15), A2 => A(15), ZN => n87);
   U62 : INV_X1 port map( A => n28, ZN => n406);
   U63 : INV_X1 port map( A => n53, ZN => n413);
   U64 : INV_X1 port map( A => n35, ZN => n409);
   U65 : INV_X1 port map( A => n52, ZN => n412);
   U66 : INV_X1 port map( A => n34, ZN => n408);
   U67 : INV_X1 port map( A => n78, ZN => n405);
   U68 : INV_X1 port map( A => n58, ZN => n411);
   U69 : INV_X1 port map( A => n39, ZN => n407);
   U70 : INV_X1 port map( A => n66, ZN => n414);
   U72 : INV_X1 port map( A => n46, ZN => n410);
   U73 : INV_X1 port map( A => n25, ZN => n415);
   U74 : NOR2_X1 port map( A1 => B(21), A2 => A(21), ZN => n52);
   U75 : NOR2_X1 port map( A1 => B(25), A2 => A(25), ZN => n34);
   U76 : NAND2_X1 port map( A1 => n87, A2 => n398, ZN => n88);
   U77 : INV_X1 port map( A => n85, ZN => n398);
   U78 : NOR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n62);
   U79 : NOR2_X1 port map( A1 => B(24), A2 => A(24), ZN => n42);
   U80 : NOR2_X1 port map( A1 => B(28), A2 => A(28), ZN => n25);
   U81 : NOR2_X1 port map( A1 => B(19), A2 => A(19), ZN => n66);
   U82 : NOR2_X1 port map( A1 => B(23), A2 => A(23), ZN => n46);
   U83 : NOR2_X1 port map( A1 => B(27), A2 => A(27), ZN => n28);
   U84 : OR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n70);
   U85 : OR2_X1 port map( A1 => B(22), A2 => A(22), ZN => n50);
   U86 : OR2_X1 port map( A1 => B(26), A2 => A(26), ZN => n32);
   U87 : NAND2_X1 port map( A1 => B(21), A2 => A(21), ZN => n54);
   U88 : NAND2_X1 port map( A1 => B(25), A2 => A(25), ZN => n36);
   U89 : NAND2_X1 port map( A1 => B(27), A2 => A(27), ZN => n29);
   U90 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n53);
   U91 : NAND2_X1 port map( A1 => B(24), A2 => A(24), ZN => n35);
   U92 : NAND2_X1 port map( A1 => B(18), A2 => A(18), ZN => n78);
   U93 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => n58);
   U94 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => n39);
   U95 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n67);
   U96 : NAND2_X1 port map( A1 => B(23), A2 => A(23), ZN => n47);
   U97 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n24);
   U98 : INV_X1 port map( A => n84, ZN => n401);
   U99 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n84);
   U101 : XNOR2_X1 port map( A => B(29), B => A(29), ZN => n21);
   U102 : AOI21_X1 port map( B1 => n23, B2 => n415, A => n24, ZN => n22);
   U103 : NAND2_X1 port map( A1 => B(14), A2 => A(14), ZN => n86);
   U104 : INV_X1 port map( A => n89, ZN => SUM_14_port);
   U105 : OAI21_X1 port map( B1 => B(14), B2 => A(14), A => n86, ZN => n89);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW02_mult_0 is

   port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  PRODUCT
         : out std_logic_vector (31 downto 0));

end ALU_N32_DW02_mult_0;

architecture SYN_csa of ALU_N32_DW02_mult_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ALU_N32_DW01_add_1_DW01_add_3
      port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (29 downto 0);  CO : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal ab_15_15_port, ab_15_14_port, ab_15_13_port, ab_15_12_port, 
      ab_15_11_port, ab_15_10_port, ab_15_9_port, ab_15_8_port, ab_15_7_port, 
      ab_15_6_port, ab_15_5_port, ab_15_4_port, ab_15_3_port, ab_15_2_port, 
      ab_15_1_port, ab_15_0_port, ab_14_15_port, ab_14_14_port, ab_14_13_port, 
      ab_14_12_port, ab_14_11_port, ab_14_10_port, ab_14_9_port, ab_14_8_port, 
      ab_14_7_port, ab_14_6_port, ab_14_5_port, ab_14_4_port, ab_14_3_port, 
      ab_14_2_port, ab_14_1_port, ab_14_0_port, ab_13_15_port, ab_13_14_port, 
      ab_13_13_port, ab_13_12_port, ab_13_11_port, ab_13_10_port, ab_13_9_port,
      ab_13_8_port, ab_13_7_port, ab_13_6_port, ab_13_5_port, ab_13_4_port, 
      ab_13_3_port, ab_13_2_port, ab_13_1_port, ab_13_0_port, ab_12_15_port, 
      ab_12_14_port, ab_12_13_port, ab_12_12_port, ab_12_11_port, ab_12_10_port
      , ab_12_9_port, ab_12_8_port, ab_12_7_port, ab_12_6_port, ab_12_5_port, 
      ab_12_4_port, ab_12_3_port, ab_12_2_port, ab_12_1_port, ab_12_0_port, 
      ab_11_15_port, ab_11_14_port, ab_11_13_port, ab_11_12_port, ab_11_11_port
      , ab_11_10_port, ab_11_9_port, ab_11_8_port, ab_11_7_port, ab_11_6_port, 
      ab_11_5_port, ab_11_4_port, ab_11_3_port, ab_11_2_port, ab_11_1_port, 
      ab_11_0_port, ab_10_15_port, ab_10_14_port, ab_10_13_port, ab_10_12_port,
      ab_10_11_port, ab_10_10_port, ab_10_9_port, ab_10_8_port, ab_10_7_port, 
      ab_10_6_port, ab_10_5_port, ab_10_4_port, ab_10_3_port, ab_10_2_port, 
      ab_10_1_port, ab_10_0_port, ab_9_15_port, ab_9_14_port, ab_9_13_port, 
      ab_9_12_port, ab_9_11_port, ab_9_10_port, ab_9_9_port, ab_9_8_port, 
      ab_9_7_port, ab_9_6_port, ab_9_5_port, ab_9_4_port, ab_9_3_port, 
      ab_9_2_port, ab_9_1_port, ab_9_0_port, ab_8_15_port, ab_8_14_port, 
      ab_8_13_port, ab_8_12_port, ab_8_11_port, ab_8_10_port, ab_8_9_port, 
      ab_8_8_port, ab_8_7_port, ab_8_6_port, ab_8_5_port, ab_8_4_port, 
      ab_8_3_port, ab_8_2_port, ab_8_1_port, ab_8_0_port, ab_7_15_port, 
      ab_7_14_port, ab_7_13_port, ab_7_12_port, ab_7_11_port, ab_7_10_port, 
      ab_7_9_port, ab_7_8_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, 
      ab_7_4_port, ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, 
      ab_6_15_port, ab_6_14_port, ab_6_13_port, ab_6_12_port, ab_6_11_port, 
      ab_6_10_port, ab_6_9_port, ab_6_8_port, ab_6_7_port, ab_6_6_port, 
      ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, ab_6_1_port, 
      ab_6_0_port, ab_5_15_port, ab_5_14_port, ab_5_13_port, ab_5_12_port, 
      ab_5_11_port, ab_5_10_port, ab_5_9_port, ab_5_8_port, ab_5_7_port, 
      ab_5_6_port, ab_5_5_port, ab_5_4_port, ab_5_3_port, ab_5_2_port, 
      ab_5_1_port, ab_5_0_port, ab_4_15_port, ab_4_14_port, ab_4_13_port, 
      ab_4_12_port, ab_4_11_port, ab_4_10_port, ab_4_9_port, ab_4_8_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_15_port, ab_3_14_port, 
      ab_3_13_port, ab_3_12_port, ab_3_11_port, ab_3_10_port, ab_3_9_port, 
      ab_3_8_port, ab_3_7_port, ab_3_6_port, ab_3_5_port, ab_3_4_port, 
      ab_3_3_port, ab_3_2_port, ab_3_1_port, ab_3_0_port, ab_2_15_port, 
      ab_2_14_port, ab_2_13_port, ab_2_12_port, ab_2_11_port, ab_2_10_port, 
      ab_2_9_port, ab_2_8_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, 
      ab_2_4_port, ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, 
      ab_1_15_port, ab_1_14_port, ab_1_13_port, ab_1_12_port, ab_1_11_port, 
      ab_1_10_port, ab_1_9_port, ab_1_8_port, ab_1_7_port, ab_1_6_port, 
      ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, ab_1_1_port, 
      ab_1_0_port, ab_0_15_port, ab_0_14_port, ab_0_13_port, ab_0_12_port, 
      ab_0_11_port, ab_0_10_port, ab_0_9_port, ab_0_8_port, ab_0_7_port, 
      ab_0_6_port, ab_0_5_port, ab_0_4_port, ab_0_3_port, ab_0_2_port, 
      ab_0_1_port, CARRYB_15_15_port, CARRYB_15_14_port, CARRYB_15_13_port, 
      CARRYB_15_12_port, CARRYB_15_11_port, CARRYB_15_10_port, CARRYB_15_9_port
      , CARRYB_15_8_port, CARRYB_15_7_port, CARRYB_15_6_port, CARRYB_15_5_port,
      CARRYB_15_4_port, CARRYB_15_3_port, CARRYB_15_2_port, CARRYB_15_1_port, 
      CARRYB_15_0_port, CARRYB_14_14_port, CARRYB_14_13_port, CARRYB_14_12_port
      , CARRYB_14_11_port, CARRYB_14_10_port, CARRYB_14_9_port, 
      CARRYB_14_8_port, CARRYB_14_7_port, CARRYB_14_6_port, CARRYB_14_5_port, 
      CARRYB_14_4_port, CARRYB_14_3_port, CARRYB_14_2_port, CARRYB_14_1_port, 
      CARRYB_14_0_port, CARRYB_13_14_port, CARRYB_13_13_port, CARRYB_13_12_port
      , CARRYB_13_11_port, CARRYB_13_10_port, CARRYB_13_9_port, 
      CARRYB_13_8_port, CARRYB_13_7_port, CARRYB_13_6_port, CARRYB_13_5_port, 
      CARRYB_13_4_port, CARRYB_13_3_port, CARRYB_13_2_port, CARRYB_13_1_port, 
      CARRYB_13_0_port, CARRYB_12_14_port, CARRYB_12_13_port, CARRYB_12_12_port
      , CARRYB_12_11_port, CARRYB_12_10_port, CARRYB_12_9_port, 
      CARRYB_12_8_port, CARRYB_12_7_port, CARRYB_12_6_port, CARRYB_12_5_port, 
      CARRYB_12_4_port, CARRYB_12_3_port, CARRYB_12_2_port, CARRYB_12_1_port, 
      CARRYB_12_0_port, CARRYB_11_14_port, CARRYB_11_13_port, CARRYB_11_12_port
      , CARRYB_11_11_port, CARRYB_11_10_port, CARRYB_11_9_port, 
      CARRYB_11_8_port, CARRYB_11_7_port, CARRYB_11_6_port, CARRYB_11_5_port, 
      CARRYB_11_4_port, CARRYB_11_3_port, CARRYB_11_2_port, CARRYB_11_1_port, 
      CARRYB_11_0_port, CARRYB_10_14_port, CARRYB_10_13_port, CARRYB_10_12_port
      , CARRYB_10_11_port, CARRYB_10_10_port, CARRYB_10_9_port, 
      CARRYB_10_8_port, CARRYB_10_7_port, CARRYB_10_6_port, CARRYB_10_5_port, 
      CARRYB_10_4_port, CARRYB_10_3_port, CARRYB_10_2_port, CARRYB_10_1_port, 
      CARRYB_10_0_port, CARRYB_9_14_port, CARRYB_9_13_port, CARRYB_9_12_port, 
      CARRYB_9_11_port, CARRYB_9_10_port, CARRYB_9_9_port, CARRYB_9_8_port, 
      CARRYB_9_7_port, CARRYB_9_6_port, CARRYB_9_5_port, CARRYB_9_4_port, 
      CARRYB_9_3_port, CARRYB_9_2_port, CARRYB_9_1_port, CARRYB_9_0_port, 
      CARRYB_8_14_port, CARRYB_8_13_port, CARRYB_8_12_port, CARRYB_8_11_port, 
      CARRYB_8_10_port, CARRYB_8_9_port, CARRYB_8_8_port, CARRYB_8_7_port, 
      CARRYB_8_6_port, CARRYB_8_5_port, CARRYB_8_4_port, CARRYB_8_3_port, 
      CARRYB_8_2_port, CARRYB_8_1_port, CARRYB_8_0_port, CARRYB_7_14_port, 
      CARRYB_7_13_port, CARRYB_7_12_port, CARRYB_7_11_port, CARRYB_7_10_port, 
      CARRYB_7_9_port, CARRYB_7_8_port, CARRYB_7_7_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_14_port, CARRYB_6_13_port, 
      CARRYB_6_12_port, CARRYB_6_11_port, CARRYB_6_10_port, CARRYB_6_9_port, 
      CARRYB_6_8_port, CARRYB_6_7_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_14_port, CARRYB_5_13_port, CARRYB_5_12_port, 
      CARRYB_5_11_port, CARRYB_5_10_port, CARRYB_5_9_port, CARRYB_5_8_port, 
      CARRYB_5_7_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_14_port, CARRYB_4_13_port, CARRYB_4_12_port, CARRYB_4_11_port, 
      CARRYB_4_10_port, CARRYB_4_9_port, CARRYB_4_8_port, CARRYB_4_7_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_14_port, 
      CARRYB_3_13_port, CARRYB_3_12_port, CARRYB_3_11_port, CARRYB_3_10_port, 
      CARRYB_3_9_port, CARRYB_3_8_port, CARRYB_3_7_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_14_port, CARRYB_2_13_port, 
      CARRYB_2_12_port, CARRYB_2_11_port, CARRYB_2_10_port, CARRYB_2_9_port, 
      CARRYB_2_8_port, CARRYB_2_7_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_15_15_port, SUMB_15_14_port, SUMB_15_13_port, 
      SUMB_15_12_port, SUMB_15_11_port, SUMB_15_10_port, SUMB_15_9_port, 
      SUMB_15_8_port, SUMB_15_7_port, SUMB_15_6_port, SUMB_15_5_port, 
      SUMB_15_4_port, SUMB_15_3_port, SUMB_15_2_port, SUMB_15_1_port, 
      SUMB_15_0_port, SUMB_14_14_port, SUMB_14_13_port, SUMB_14_12_port, 
      SUMB_14_11_port, SUMB_14_10_port, SUMB_14_9_port, SUMB_14_8_port, 
      SUMB_14_7_port, SUMB_14_6_port, SUMB_14_5_port, SUMB_14_4_port, 
      SUMB_14_3_port, SUMB_14_2_port, SUMB_14_1_port, SUMB_13_14_port, 
      SUMB_13_13_port, SUMB_13_12_port, SUMB_13_11_port, SUMB_13_10_port, 
      SUMB_13_9_port, SUMB_13_8_port, SUMB_13_7_port, SUMB_13_6_port, 
      SUMB_13_5_port, SUMB_13_4_port, SUMB_13_3_port, SUMB_13_2_port, 
      SUMB_13_1_port, SUMB_12_14_port, SUMB_12_13_port, SUMB_12_12_port, 
      SUMB_12_11_port, SUMB_12_10_port, SUMB_12_9_port, SUMB_12_8_port, 
      SUMB_12_7_port, SUMB_12_6_port, SUMB_12_5_port, SUMB_12_4_port, 
      SUMB_12_3_port, SUMB_12_2_port, SUMB_12_1_port, SUMB_11_14_port, 
      SUMB_11_13_port, SUMB_11_12_port, SUMB_11_11_port, SUMB_11_10_port, 
      SUMB_11_9_port, SUMB_11_8_port, SUMB_11_7_port, SUMB_11_6_port, 
      SUMB_11_5_port, SUMB_11_4_port, SUMB_11_3_port, SUMB_11_2_port, 
      SUMB_11_1_port, SUMB_10_14_port, SUMB_10_13_port, SUMB_10_12_port, 
      SUMB_10_11_port, SUMB_10_10_port, SUMB_10_9_port, SUMB_10_8_port, 
      SUMB_10_7_port, SUMB_10_6_port, SUMB_10_5_port, SUMB_10_4_port, 
      SUMB_10_3_port, SUMB_10_2_port, SUMB_10_1_port, SUMB_9_14_port, 
      SUMB_9_13_port, SUMB_9_12_port, SUMB_9_11_port, SUMB_9_10_port, 
      SUMB_9_9_port, SUMB_9_8_port, SUMB_9_7_port, SUMB_9_6_port, SUMB_9_5_port
      , SUMB_9_4_port, SUMB_9_3_port, SUMB_9_2_port, SUMB_9_1_port, 
      SUMB_8_14_port, SUMB_8_13_port, SUMB_8_12_port, SUMB_8_11_port, 
      SUMB_8_10_port, SUMB_8_9_port, SUMB_8_8_port, SUMB_8_7_port, 
      SUMB_8_6_port, SUMB_8_5_port, SUMB_8_4_port, SUMB_8_3_port, SUMB_8_2_port
      , SUMB_8_1_port, SUMB_7_14_port, SUMB_7_13_port, SUMB_7_12_port, 
      SUMB_7_11_port, SUMB_7_10_port, SUMB_7_9_port, SUMB_7_8_port, 
      SUMB_7_7_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, SUMB_7_3_port
      , SUMB_7_2_port, SUMB_7_1_port, SUMB_6_14_port, SUMB_6_13_port, 
      SUMB_6_12_port, SUMB_6_11_port, SUMB_6_10_port, SUMB_6_9_port, 
      SUMB_6_8_port, SUMB_6_7_port, SUMB_6_6_port, SUMB_6_5_port, SUMB_6_4_port
      , SUMB_6_3_port, SUMB_6_2_port, SUMB_6_1_port, SUMB_5_14_port, 
      SUMB_5_13_port, SUMB_5_12_port, SUMB_5_11_port, SUMB_5_10_port, 
      SUMB_5_9_port, SUMB_5_8_port, SUMB_5_7_port, SUMB_5_6_port, SUMB_5_5_port
      , SUMB_5_4_port, SUMB_5_3_port, SUMB_5_2_port, SUMB_5_1_port, 
      SUMB_4_14_port, SUMB_4_13_port, SUMB_4_12_port, SUMB_4_11_port, 
      SUMB_4_10_port, SUMB_4_9_port, SUMB_4_8_port, SUMB_4_7_port, 
      SUMB_4_6_port, SUMB_4_5_port, SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port
      , SUMB_4_1_port, SUMB_3_14_port, SUMB_3_13_port, SUMB_3_12_port, 
      SUMB_3_11_port, SUMB_3_10_port, SUMB_3_9_port, SUMB_3_8_port, 
      SUMB_3_7_port, SUMB_3_6_port, SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port
      , SUMB_3_2_port, SUMB_3_1_port, SUMB_2_14_port, SUMB_2_13_port, 
      SUMB_2_12_port, SUMB_2_11_port, SUMB_2_10_port, SUMB_2_9_port, 
      SUMB_2_8_port, SUMB_2_7_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port
      , SUMB_2_3_port, SUMB_2_2_port, SUMB_2_1_port, A1_13_port, A1_12_port, 
      A1_11_port, A1_10_port, A1_9_port, A1_8_port, A1_7_port, A1_6_port, 
      A1_5_port, A1_4_port, A1_3_port, A1_2_port, A1_1_port, A1_0_port, 
      A2_14_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n_1017 : std_logic;

begin
   
   S14_15_0 : FA_X1 port map( A => A(15), B => B(15), CI => SUMB_15_0_port, CO 
                           => A2_14_port, S => A1_13_port);
   S4_0 : FA_X1 port map( A => ab_15_0_port, B => CARRYB_14_0_port, CI => 
                           SUMB_14_1_port, CO => CARRYB_15_0_port, S => 
                           SUMB_15_0_port);
   S4_1 : FA_X1 port map( A => ab_15_1_port, B => CARRYB_14_1_port, CI => 
                           SUMB_14_2_port, CO => CARRYB_15_1_port, S => 
                           SUMB_15_1_port);
   S4_2 : FA_X1 port map( A => ab_15_2_port, B => CARRYB_14_2_port, CI => 
                           SUMB_14_3_port, CO => CARRYB_15_2_port, S => 
                           SUMB_15_2_port);
   S4_3 : FA_X1 port map( A => ab_15_3_port, B => CARRYB_14_3_port, CI => 
                           SUMB_14_4_port, CO => CARRYB_15_3_port, S => 
                           SUMB_15_3_port);
   S4_4 : FA_X1 port map( A => ab_15_4_port, B => CARRYB_14_4_port, CI => 
                           SUMB_14_5_port, CO => CARRYB_15_4_port, S => 
                           SUMB_15_4_port);
   S4_5 : FA_X1 port map( A => ab_15_5_port, B => CARRYB_14_5_port, CI => 
                           SUMB_14_6_port, CO => CARRYB_15_5_port, S => 
                           SUMB_15_5_port);
   S4_6 : FA_X1 port map( A => ab_15_6_port, B => CARRYB_14_6_port, CI => 
                           SUMB_14_7_port, CO => CARRYB_15_6_port, S => 
                           SUMB_15_6_port);
   S4_7 : FA_X1 port map( A => ab_15_7_port, B => CARRYB_14_7_port, CI => 
                           SUMB_14_8_port, CO => CARRYB_15_7_port, S => 
                           SUMB_15_7_port);
   S4_8 : FA_X1 port map( A => ab_15_8_port, B => CARRYB_14_8_port, CI => 
                           SUMB_14_9_port, CO => CARRYB_15_8_port, S => 
                           SUMB_15_8_port);
   S4_9 : FA_X1 port map( A => ab_15_9_port, B => CARRYB_14_9_port, CI => 
                           SUMB_14_10_port, CO => CARRYB_15_9_port, S => 
                           SUMB_15_9_port);
   S4_10 : FA_X1 port map( A => ab_15_10_port, B => CARRYB_14_10_port, CI => 
                           SUMB_14_11_port, CO => CARRYB_15_10_port, S => 
                           SUMB_15_10_port);
   S4_11 : FA_X1 port map( A => ab_15_11_port, B => CARRYB_14_11_port, CI => 
                           SUMB_14_12_port, CO => CARRYB_15_11_port, S => 
                           SUMB_15_11_port);
   S4_12 : FA_X1 port map( A => ab_15_12_port, B => CARRYB_14_12_port, CI => 
                           SUMB_14_13_port, CO => CARRYB_15_12_port, S => 
                           SUMB_15_12_port);
   S4_13 : FA_X1 port map( A => ab_15_13_port, B => CARRYB_14_13_port, CI => 
                           SUMB_14_14_port, CO => CARRYB_15_13_port, S => 
                           SUMB_15_13_port);
   S5_14 : FA_X1 port map( A => ab_15_14_port, B => CARRYB_14_14_port, CI => 
                           ab_14_15_port, CO => CARRYB_15_14_port, S => 
                           SUMB_15_14_port);
   S14_15 : FA_X1 port map( A => n809, B => n820, CI => ab_15_15_port, CO => 
                           CARRYB_15_15_port, S => SUMB_15_15_port);
   S1_14_0 : FA_X1 port map( A => ab_14_0_port, B => CARRYB_13_0_port, CI => 
                           SUMB_13_1_port, CO => CARRYB_14_0_port, S => 
                           A1_12_port);
   S2_14_1 : FA_X1 port map( A => ab_14_1_port, B => CARRYB_13_1_port, CI => 
                           SUMB_13_2_port, CO => CARRYB_14_1_port, S => 
                           SUMB_14_1_port);
   S2_14_2 : FA_X1 port map( A => ab_14_2_port, B => CARRYB_13_2_port, CI => 
                           SUMB_13_3_port, CO => CARRYB_14_2_port, S => 
                           SUMB_14_2_port);
   S2_14_3 : FA_X1 port map( A => ab_14_3_port, B => CARRYB_13_3_port, CI => 
                           SUMB_13_4_port, CO => CARRYB_14_3_port, S => 
                           SUMB_14_3_port);
   S2_14_4 : FA_X1 port map( A => ab_14_4_port, B => CARRYB_13_4_port, CI => 
                           SUMB_13_5_port, CO => CARRYB_14_4_port, S => 
                           SUMB_14_4_port);
   S2_14_5 : FA_X1 port map( A => ab_14_5_port, B => CARRYB_13_5_port, CI => 
                           SUMB_13_6_port, CO => CARRYB_14_5_port, S => 
                           SUMB_14_5_port);
   S2_14_6 : FA_X1 port map( A => ab_14_6_port, B => CARRYB_13_6_port, CI => 
                           SUMB_13_7_port, CO => CARRYB_14_6_port, S => 
                           SUMB_14_6_port);
   S2_14_7 : FA_X1 port map( A => ab_14_7_port, B => CARRYB_13_7_port, CI => 
                           SUMB_13_8_port, CO => CARRYB_14_7_port, S => 
                           SUMB_14_7_port);
   S2_14_8 : FA_X1 port map( A => ab_14_8_port, B => CARRYB_13_8_port, CI => 
                           SUMB_13_9_port, CO => CARRYB_14_8_port, S => 
                           SUMB_14_8_port);
   S2_14_9 : FA_X1 port map( A => ab_14_9_port, B => CARRYB_13_9_port, CI => 
                           SUMB_13_10_port, CO => CARRYB_14_9_port, S => 
                           SUMB_14_9_port);
   S2_14_10 : FA_X1 port map( A => ab_14_10_port, B => CARRYB_13_10_port, CI =>
                           SUMB_13_11_port, CO => CARRYB_14_10_port, S => 
                           SUMB_14_10_port);
   S2_14_11 : FA_X1 port map( A => ab_14_11_port, B => CARRYB_13_11_port, CI =>
                           SUMB_13_12_port, CO => CARRYB_14_11_port, S => 
                           SUMB_14_11_port);
   S2_14_12 : FA_X1 port map( A => ab_14_12_port, B => CARRYB_13_12_port, CI =>
                           SUMB_13_13_port, CO => CARRYB_14_12_port, S => 
                           SUMB_14_12_port);
   S2_14_13 : FA_X1 port map( A => ab_14_13_port, B => CARRYB_13_13_port, CI =>
                           SUMB_13_14_port, CO => CARRYB_14_13_port, S => 
                           SUMB_14_13_port);
   S3_14_14 : FA_X1 port map( A => ab_14_14_port, B => CARRYB_13_14_port, CI =>
                           ab_13_15_port, CO => CARRYB_14_14_port, S => 
                           SUMB_14_14_port);
   S1_13_0 : FA_X1 port map( A => ab_13_0_port, B => CARRYB_12_0_port, CI => 
                           SUMB_12_1_port, CO => CARRYB_13_0_port, S => 
                           A1_11_port);
   S2_13_1 : FA_X1 port map( A => ab_13_1_port, B => CARRYB_12_1_port, CI => 
                           SUMB_12_2_port, CO => CARRYB_13_1_port, S => 
                           SUMB_13_1_port);
   S2_13_2 : FA_X1 port map( A => ab_13_2_port, B => CARRYB_12_2_port, CI => 
                           SUMB_12_3_port, CO => CARRYB_13_2_port, S => 
                           SUMB_13_2_port);
   S2_13_3 : FA_X1 port map( A => ab_13_3_port, B => CARRYB_12_3_port, CI => 
                           SUMB_12_4_port, CO => CARRYB_13_3_port, S => 
                           SUMB_13_3_port);
   S2_13_4 : FA_X1 port map( A => ab_13_4_port, B => CARRYB_12_4_port, CI => 
                           SUMB_12_5_port, CO => CARRYB_13_4_port, S => 
                           SUMB_13_4_port);
   S2_13_5 : FA_X1 port map( A => ab_13_5_port, B => CARRYB_12_5_port, CI => 
                           SUMB_12_6_port, CO => CARRYB_13_5_port, S => 
                           SUMB_13_5_port);
   S2_13_6 : FA_X1 port map( A => ab_13_6_port, B => CARRYB_12_6_port, CI => 
                           SUMB_12_7_port, CO => CARRYB_13_6_port, S => 
                           SUMB_13_6_port);
   S2_13_7 : FA_X1 port map( A => ab_13_7_port, B => CARRYB_12_7_port, CI => 
                           SUMB_12_8_port, CO => CARRYB_13_7_port, S => 
                           SUMB_13_7_port);
   S2_13_8 : FA_X1 port map( A => ab_13_8_port, B => CARRYB_12_8_port, CI => 
                           SUMB_12_9_port, CO => CARRYB_13_8_port, S => 
                           SUMB_13_8_port);
   S2_13_9 : FA_X1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, CI => 
                           SUMB_12_10_port, CO => CARRYB_13_9_port, S => 
                           SUMB_13_9_port);
   S2_13_10 : FA_X1 port map( A => ab_13_10_port, B => CARRYB_12_10_port, CI =>
                           SUMB_12_11_port, CO => CARRYB_13_10_port, S => 
                           SUMB_13_10_port);
   S2_13_11 : FA_X1 port map( A => ab_13_11_port, B => CARRYB_12_11_port, CI =>
                           SUMB_12_12_port, CO => CARRYB_13_11_port, S => 
                           SUMB_13_11_port);
   S2_13_12 : FA_X1 port map( A => ab_13_12_port, B => CARRYB_12_12_port, CI =>
                           SUMB_12_13_port, CO => CARRYB_13_12_port, S => 
                           SUMB_13_12_port);
   S2_13_13 : FA_X1 port map( A => ab_13_13_port, B => CARRYB_12_13_port, CI =>
                           SUMB_12_14_port, CO => CARRYB_13_13_port, S => 
                           SUMB_13_13_port);
   S3_13_14 : FA_X1 port map( A => ab_13_14_port, B => CARRYB_12_14_port, CI =>
                           ab_12_15_port, CO => CARRYB_13_14_port, S => 
                           SUMB_13_14_port);
   S1_12_0 : FA_X1 port map( A => ab_12_0_port, B => CARRYB_11_0_port, CI => 
                           SUMB_11_1_port, CO => CARRYB_12_0_port, S => 
                           A1_10_port);
   S2_12_1 : FA_X1 port map( A => ab_12_1_port, B => CARRYB_11_1_port, CI => 
                           SUMB_11_2_port, CO => CARRYB_12_1_port, S => 
                           SUMB_12_1_port);
   S2_12_2 : FA_X1 port map( A => ab_12_2_port, B => CARRYB_11_2_port, CI => 
                           SUMB_11_3_port, CO => CARRYB_12_2_port, S => 
                           SUMB_12_2_port);
   S2_12_3 : FA_X1 port map( A => ab_12_3_port, B => CARRYB_11_3_port, CI => 
                           SUMB_11_4_port, CO => CARRYB_12_3_port, S => 
                           SUMB_12_3_port);
   S2_12_4 : FA_X1 port map( A => ab_12_4_port, B => CARRYB_11_4_port, CI => 
                           SUMB_11_5_port, CO => CARRYB_12_4_port, S => 
                           SUMB_12_4_port);
   S2_12_5 : FA_X1 port map( A => ab_12_5_port, B => CARRYB_11_5_port, CI => 
                           SUMB_11_6_port, CO => CARRYB_12_5_port, S => 
                           SUMB_12_5_port);
   S2_12_6 : FA_X1 port map( A => ab_12_6_port, B => CARRYB_11_6_port, CI => 
                           SUMB_11_7_port, CO => CARRYB_12_6_port, S => 
                           SUMB_12_6_port);
   S2_12_7 : FA_X1 port map( A => ab_12_7_port, B => CARRYB_11_7_port, CI => 
                           SUMB_11_8_port, CO => CARRYB_12_7_port, S => 
                           SUMB_12_7_port);
   S2_12_8 : FA_X1 port map( A => ab_12_8_port, B => CARRYB_11_8_port, CI => 
                           SUMB_11_9_port, CO => CARRYB_12_8_port, S => 
                           SUMB_12_8_port);
   S2_12_9 : FA_X1 port map( A => ab_12_9_port, B => CARRYB_11_9_port, CI => 
                           SUMB_11_10_port, CO => CARRYB_12_9_port, S => 
                           SUMB_12_9_port);
   S2_12_10 : FA_X1 port map( A => ab_12_10_port, B => CARRYB_11_10_port, CI =>
                           SUMB_11_11_port, CO => CARRYB_12_10_port, S => 
                           SUMB_12_10_port);
   S2_12_11 : FA_X1 port map( A => ab_12_11_port, B => CARRYB_11_11_port, CI =>
                           SUMB_11_12_port, CO => CARRYB_12_11_port, S => 
                           SUMB_12_11_port);
   S2_12_12 : FA_X1 port map( A => ab_12_12_port, B => CARRYB_11_12_port, CI =>
                           SUMB_11_13_port, CO => CARRYB_12_12_port, S => 
                           SUMB_12_12_port);
   S2_12_13 : FA_X1 port map( A => ab_12_13_port, B => CARRYB_11_13_port, CI =>
                           SUMB_11_14_port, CO => CARRYB_12_13_port, S => 
                           SUMB_12_13_port);
   S3_12_14 : FA_X1 port map( A => ab_12_14_port, B => CARRYB_11_14_port, CI =>
                           ab_11_15_port, CO => CARRYB_12_14_port, S => 
                           SUMB_12_14_port);
   S1_11_0 : FA_X1 port map( A => ab_11_0_port, B => CARRYB_10_0_port, CI => 
                           SUMB_10_1_port, CO => CARRYB_11_0_port, S => 
                           A1_9_port);
   S2_11_1 : FA_X1 port map( A => ab_11_1_port, B => CARRYB_10_1_port, CI => 
                           SUMB_10_2_port, CO => CARRYB_11_1_port, S => 
                           SUMB_11_1_port);
   S2_11_2 : FA_X1 port map( A => ab_11_2_port, B => CARRYB_10_2_port, CI => 
                           SUMB_10_3_port, CO => CARRYB_11_2_port, S => 
                           SUMB_11_2_port);
   S2_11_3 : FA_X1 port map( A => ab_11_3_port, B => CARRYB_10_3_port, CI => 
                           SUMB_10_4_port, CO => CARRYB_11_3_port, S => 
                           SUMB_11_3_port);
   S2_11_4 : FA_X1 port map( A => ab_11_4_port, B => CARRYB_10_4_port, CI => 
                           SUMB_10_5_port, CO => CARRYB_11_4_port, S => 
                           SUMB_11_4_port);
   S2_11_5 : FA_X1 port map( A => ab_11_5_port, B => CARRYB_10_5_port, CI => 
                           SUMB_10_6_port, CO => CARRYB_11_5_port, S => 
                           SUMB_11_5_port);
   S2_11_6 : FA_X1 port map( A => ab_11_6_port, B => CARRYB_10_6_port, CI => 
                           SUMB_10_7_port, CO => CARRYB_11_6_port, S => 
                           SUMB_11_6_port);
   S2_11_7 : FA_X1 port map( A => ab_11_7_port, B => CARRYB_10_7_port, CI => 
                           SUMB_10_8_port, CO => CARRYB_11_7_port, S => 
                           SUMB_11_7_port);
   S2_11_8 : FA_X1 port map( A => ab_11_8_port, B => CARRYB_10_8_port, CI => 
                           SUMB_10_9_port, CO => CARRYB_11_8_port, S => 
                           SUMB_11_8_port);
   S2_11_9 : FA_X1 port map( A => ab_11_9_port, B => CARRYB_10_9_port, CI => 
                           SUMB_10_10_port, CO => CARRYB_11_9_port, S => 
                           SUMB_11_9_port);
   S2_11_10 : FA_X1 port map( A => ab_11_10_port, B => CARRYB_10_10_port, CI =>
                           SUMB_10_11_port, CO => CARRYB_11_10_port, S => 
                           SUMB_11_10_port);
   S2_11_11 : FA_X1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, CI =>
                           SUMB_10_12_port, CO => CARRYB_11_11_port, S => 
                           SUMB_11_11_port);
   S2_11_12 : FA_X1 port map( A => ab_11_12_port, B => CARRYB_10_12_port, CI =>
                           SUMB_10_13_port, CO => CARRYB_11_12_port, S => 
                           SUMB_11_12_port);
   S2_11_13 : FA_X1 port map( A => ab_11_13_port, B => CARRYB_10_13_port, CI =>
                           SUMB_10_14_port, CO => CARRYB_11_13_port, S => 
                           SUMB_11_13_port);
   S3_11_14 : FA_X1 port map( A => ab_11_14_port, B => CARRYB_10_14_port, CI =>
                           ab_10_15_port, CO => CARRYB_11_14_port, S => 
                           SUMB_11_14_port);
   S1_10_0 : FA_X1 port map( A => ab_10_0_port, B => CARRYB_9_0_port, CI => 
                           SUMB_9_1_port, CO => CARRYB_10_0_port, S => 
                           A1_8_port);
   S2_10_1 : FA_X1 port map( A => ab_10_1_port, B => CARRYB_9_1_port, CI => 
                           SUMB_9_2_port, CO => CARRYB_10_1_port, S => 
                           SUMB_10_1_port);
   S2_10_2 : FA_X1 port map( A => ab_10_2_port, B => CARRYB_9_2_port, CI => 
                           SUMB_9_3_port, CO => CARRYB_10_2_port, S => 
                           SUMB_10_2_port);
   S2_10_3 : FA_X1 port map( A => ab_10_3_port, B => CARRYB_9_3_port, CI => 
                           SUMB_9_4_port, CO => CARRYB_10_3_port, S => 
                           SUMB_10_3_port);
   S2_10_4 : FA_X1 port map( A => ab_10_4_port, B => CARRYB_9_4_port, CI => 
                           SUMB_9_5_port, CO => CARRYB_10_4_port, S => 
                           SUMB_10_4_port);
   S2_10_5 : FA_X1 port map( A => ab_10_5_port, B => CARRYB_9_5_port, CI => 
                           SUMB_9_6_port, CO => CARRYB_10_5_port, S => 
                           SUMB_10_5_port);
   S2_10_6 : FA_X1 port map( A => ab_10_6_port, B => CARRYB_9_6_port, CI => 
                           SUMB_9_7_port, CO => CARRYB_10_6_port, S => 
                           SUMB_10_6_port);
   S2_10_7 : FA_X1 port map( A => ab_10_7_port, B => CARRYB_9_7_port, CI => 
                           SUMB_9_8_port, CO => CARRYB_10_7_port, S => 
                           SUMB_10_7_port);
   S2_10_8 : FA_X1 port map( A => ab_10_8_port, B => CARRYB_9_8_port, CI => 
                           SUMB_9_9_port, CO => CARRYB_10_8_port, S => 
                           SUMB_10_8_port);
   S2_10_9 : FA_X1 port map( A => ab_10_9_port, B => CARRYB_9_9_port, CI => 
                           SUMB_9_10_port, CO => CARRYB_10_9_port, S => 
                           SUMB_10_9_port);
   S2_10_10 : FA_X1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, CI => 
                           SUMB_9_11_port, CO => CARRYB_10_10_port, S => 
                           SUMB_10_10_port);
   S2_10_11 : FA_X1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, CI => 
                           SUMB_9_12_port, CO => CARRYB_10_11_port, S => 
                           SUMB_10_11_port);
   S2_10_12 : FA_X1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, CI => 
                           SUMB_9_13_port, CO => CARRYB_10_12_port, S => 
                           SUMB_10_12_port);
   S2_10_13 : FA_X1 port map( A => ab_10_13_port, B => CARRYB_9_13_port, CI => 
                           SUMB_9_14_port, CO => CARRYB_10_13_port, S => 
                           SUMB_10_13_port);
   S3_10_14 : FA_X1 port map( A => ab_10_14_port, B => CARRYB_9_14_port, CI => 
                           ab_9_15_port, CO => CARRYB_10_14_port, S => 
                           SUMB_10_14_port);
   S1_9_0 : FA_X1 port map( A => ab_9_0_port, B => CARRYB_8_0_port, CI => 
                           SUMB_8_1_port, CO => CARRYB_9_0_port, S => A1_7_port
                           );
   S2_9_1 : FA_X1 port map( A => ab_9_1_port, B => CARRYB_8_1_port, CI => 
                           SUMB_8_2_port, CO => CARRYB_9_1_port, S => 
                           SUMB_9_1_port);
   S2_9_2 : FA_X1 port map( A => ab_9_2_port, B => CARRYB_8_2_port, CI => 
                           SUMB_8_3_port, CO => CARRYB_9_2_port, S => 
                           SUMB_9_2_port);
   S2_9_3 : FA_X1 port map( A => ab_9_3_port, B => CARRYB_8_3_port, CI => 
                           SUMB_8_4_port, CO => CARRYB_9_3_port, S => 
                           SUMB_9_3_port);
   S2_9_4 : FA_X1 port map( A => ab_9_4_port, B => CARRYB_8_4_port, CI => 
                           SUMB_8_5_port, CO => CARRYB_9_4_port, S => 
                           SUMB_9_4_port);
   S2_9_5 : FA_X1 port map( A => ab_9_5_port, B => CARRYB_8_5_port, CI => 
                           SUMB_8_6_port, CO => CARRYB_9_5_port, S => 
                           SUMB_9_5_port);
   S2_9_6 : FA_X1 port map( A => ab_9_6_port, B => CARRYB_8_6_port, CI => 
                           SUMB_8_7_port, CO => CARRYB_9_6_port, S => 
                           SUMB_9_6_port);
   S2_9_7 : FA_X1 port map( A => ab_9_7_port, B => CARRYB_8_7_port, CI => 
                           SUMB_8_8_port, CO => CARRYB_9_7_port, S => 
                           SUMB_9_7_port);
   S2_9_8 : FA_X1 port map( A => ab_9_8_port, B => CARRYB_8_8_port, CI => 
                           SUMB_8_9_port, CO => CARRYB_9_8_port, S => 
                           SUMB_9_8_port);
   S2_9_9 : FA_X1 port map( A => ab_9_9_port, B => CARRYB_8_9_port, CI => 
                           SUMB_8_10_port, CO => CARRYB_9_9_port, S => 
                           SUMB_9_9_port);
   S2_9_10 : FA_X1 port map( A => ab_9_10_port, B => CARRYB_8_10_port, CI => 
                           SUMB_8_11_port, CO => CARRYB_9_10_port, S => 
                           SUMB_9_10_port);
   S2_9_11 : FA_X1 port map( A => ab_9_11_port, B => CARRYB_8_11_port, CI => 
                           SUMB_8_12_port, CO => CARRYB_9_11_port, S => 
                           SUMB_9_11_port);
   S2_9_12 : FA_X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, CI => 
                           SUMB_8_13_port, CO => CARRYB_9_12_port, S => 
                           SUMB_9_12_port);
   S2_9_13 : FA_X1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, CI => 
                           SUMB_8_14_port, CO => CARRYB_9_13_port, S => 
                           SUMB_9_13_port);
   S3_9_14 : FA_X1 port map( A => ab_9_14_port, B => CARRYB_8_14_port, CI => 
                           ab_8_15_port, CO => CARRYB_9_14_port, S => 
                           SUMB_9_14_port);
   S1_8_0 : FA_X1 port map( A => ab_8_0_port, B => CARRYB_7_0_port, CI => 
                           SUMB_7_1_port, CO => CARRYB_8_0_port, S => A1_6_port
                           );
   S2_8_1 : FA_X1 port map( A => ab_8_1_port, B => CARRYB_7_1_port, CI => 
                           SUMB_7_2_port, CO => CARRYB_8_1_port, S => 
                           SUMB_8_1_port);
   S2_8_2 : FA_X1 port map( A => ab_8_2_port, B => CARRYB_7_2_port, CI => 
                           SUMB_7_3_port, CO => CARRYB_8_2_port, S => 
                           SUMB_8_2_port);
   S2_8_3 : FA_X1 port map( A => ab_8_3_port, B => CARRYB_7_3_port, CI => 
                           SUMB_7_4_port, CO => CARRYB_8_3_port, S => 
                           SUMB_8_3_port);
   S2_8_4 : FA_X1 port map( A => ab_8_4_port, B => CARRYB_7_4_port, CI => 
                           SUMB_7_5_port, CO => CARRYB_8_4_port, S => 
                           SUMB_8_4_port);
   S2_8_5 : FA_X1 port map( A => ab_8_5_port, B => CARRYB_7_5_port, CI => 
                           SUMB_7_6_port, CO => CARRYB_8_5_port, S => 
                           SUMB_8_5_port);
   S2_8_6 : FA_X1 port map( A => ab_8_6_port, B => CARRYB_7_6_port, CI => 
                           SUMB_7_7_port, CO => CARRYB_8_6_port, S => 
                           SUMB_8_6_port);
   S2_8_7 : FA_X1 port map( A => ab_8_7_port, B => CARRYB_7_7_port, CI => 
                           SUMB_7_8_port, CO => CARRYB_8_7_port, S => 
                           SUMB_8_7_port);
   S2_8_8 : FA_X1 port map( A => ab_8_8_port, B => CARRYB_7_8_port, CI => 
                           SUMB_7_9_port, CO => CARRYB_8_8_port, S => 
                           SUMB_8_8_port);
   S2_8_9 : FA_X1 port map( A => ab_8_9_port, B => CARRYB_7_9_port, CI => 
                           SUMB_7_10_port, CO => CARRYB_8_9_port, S => 
                           SUMB_8_9_port);
   S2_8_10 : FA_X1 port map( A => ab_8_10_port, B => CARRYB_7_10_port, CI => 
                           SUMB_7_11_port, CO => CARRYB_8_10_port, S => 
                           SUMB_8_10_port);
   S2_8_11 : FA_X1 port map( A => ab_8_11_port, B => CARRYB_7_11_port, CI => 
                           SUMB_7_12_port, CO => CARRYB_8_11_port, S => 
                           SUMB_8_11_port);
   S2_8_12 : FA_X1 port map( A => ab_8_12_port, B => CARRYB_7_12_port, CI => 
                           SUMB_7_13_port, CO => CARRYB_8_12_port, S => 
                           SUMB_8_12_port);
   S2_8_13 : FA_X1 port map( A => ab_8_13_port, B => CARRYB_7_13_port, CI => 
                           SUMB_7_14_port, CO => CARRYB_8_13_port, S => 
                           SUMB_8_13_port);
   S3_8_14 : FA_X1 port map( A => ab_8_14_port, B => CARRYB_7_14_port, CI => 
                           ab_7_15_port, CO => CARRYB_8_14_port, S => 
                           SUMB_8_14_port);
   S1_7_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => A1_5_port
                           );
   S2_7_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S2_7_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S2_7_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S2_7_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S2_7_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S2_7_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           SUMB_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S2_7_7 : FA_X1 port map( A => ab_7_7_port, B => CARRYB_6_7_port, CI => 
                           SUMB_6_8_port, CO => CARRYB_7_7_port, S => 
                           SUMB_7_7_port);
   S2_7_8 : FA_X1 port map( A => ab_7_8_port, B => CARRYB_6_8_port, CI => 
                           SUMB_6_9_port, CO => CARRYB_7_8_port, S => 
                           SUMB_7_8_port);
   S2_7_9 : FA_X1 port map( A => ab_7_9_port, B => CARRYB_6_9_port, CI => 
                           SUMB_6_10_port, CO => CARRYB_7_9_port, S => 
                           SUMB_7_9_port);
   S2_7_10 : FA_X1 port map( A => ab_7_10_port, B => CARRYB_6_10_port, CI => 
                           SUMB_6_11_port, CO => CARRYB_7_10_port, S => 
                           SUMB_7_10_port);
   S2_7_11 : FA_X1 port map( A => ab_7_11_port, B => CARRYB_6_11_port, CI => 
                           SUMB_6_12_port, CO => CARRYB_7_11_port, S => 
                           SUMB_7_11_port);
   S2_7_12 : FA_X1 port map( A => ab_7_12_port, B => CARRYB_6_12_port, CI => 
                           SUMB_6_13_port, CO => CARRYB_7_12_port, S => 
                           SUMB_7_12_port);
   S2_7_13 : FA_X1 port map( A => ab_7_13_port, B => CARRYB_6_13_port, CI => 
                           SUMB_6_14_port, CO => CARRYB_7_13_port, S => 
                           SUMB_7_13_port);
   S3_7_14 : FA_X1 port map( A => ab_7_14_port, B => CARRYB_6_14_port, CI => 
                           ab_6_15_port, CO => CARRYB_7_14_port, S => 
                           SUMB_7_14_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S2_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           SUMB_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S2_6_7 : FA_X1 port map( A => ab_6_7_port, B => CARRYB_5_7_port, CI => 
                           SUMB_5_8_port, CO => CARRYB_6_7_port, S => 
                           SUMB_6_7_port);
   S2_6_8 : FA_X1 port map( A => ab_6_8_port, B => CARRYB_5_8_port, CI => 
                           SUMB_5_9_port, CO => CARRYB_6_8_port, S => 
                           SUMB_6_8_port);
   S2_6_9 : FA_X1 port map( A => ab_6_9_port, B => CARRYB_5_9_port, CI => 
                           SUMB_5_10_port, CO => CARRYB_6_9_port, S => 
                           SUMB_6_9_port);
   S2_6_10 : FA_X1 port map( A => ab_6_10_port, B => CARRYB_5_10_port, CI => 
                           SUMB_5_11_port, CO => CARRYB_6_10_port, S => 
                           SUMB_6_10_port);
   S2_6_11 : FA_X1 port map( A => ab_6_11_port, B => CARRYB_5_11_port, CI => 
                           SUMB_5_12_port, CO => CARRYB_6_11_port, S => 
                           SUMB_6_11_port);
   S2_6_12 : FA_X1 port map( A => ab_6_12_port, B => CARRYB_5_12_port, CI => 
                           SUMB_5_13_port, CO => CARRYB_6_12_port, S => 
                           SUMB_6_12_port);
   S2_6_13 : FA_X1 port map( A => ab_6_13_port, B => CARRYB_5_13_port, CI => 
                           SUMB_5_14_port, CO => CARRYB_6_13_port, S => 
                           SUMB_6_13_port);
   S3_6_14 : FA_X1 port map( A => ab_6_14_port, B => CARRYB_5_14_port, CI => 
                           ab_5_15_port, CO => CARRYB_6_14_port, S => 
                           SUMB_6_14_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S2_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           SUMB_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S2_5_7 : FA_X1 port map( A => ab_5_7_port, B => CARRYB_4_7_port, CI => 
                           SUMB_4_8_port, CO => CARRYB_5_7_port, S => 
                           SUMB_5_7_port);
   S2_5_8 : FA_X1 port map( A => ab_5_8_port, B => CARRYB_4_8_port, CI => 
                           SUMB_4_9_port, CO => CARRYB_5_8_port, S => 
                           SUMB_5_8_port);
   S2_5_9 : FA_X1 port map( A => ab_5_9_port, B => CARRYB_4_9_port, CI => 
                           SUMB_4_10_port, CO => CARRYB_5_9_port, S => 
                           SUMB_5_9_port);
   S2_5_10 : FA_X1 port map( A => ab_5_10_port, B => CARRYB_4_10_port, CI => 
                           SUMB_4_11_port, CO => CARRYB_5_10_port, S => 
                           SUMB_5_10_port);
   S2_5_11 : FA_X1 port map( A => ab_5_11_port, B => CARRYB_4_11_port, CI => 
                           SUMB_4_12_port, CO => CARRYB_5_11_port, S => 
                           SUMB_5_11_port);
   S2_5_12 : FA_X1 port map( A => ab_5_12_port, B => CARRYB_4_12_port, CI => 
                           SUMB_4_13_port, CO => CARRYB_5_12_port, S => 
                           SUMB_5_12_port);
   S2_5_13 : FA_X1 port map( A => ab_5_13_port, B => CARRYB_4_13_port, CI => 
                           SUMB_4_14_port, CO => CARRYB_5_13_port, S => 
                           SUMB_5_13_port);
   S3_5_14 : FA_X1 port map( A => ab_5_14_port, B => CARRYB_4_14_port, CI => 
                           ab_4_15_port, CO => CARRYB_5_14_port, S => 
                           SUMB_5_14_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S2_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           SUMB_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S2_4_7 : FA_X1 port map( A => ab_4_7_port, B => CARRYB_3_7_port, CI => 
                           SUMB_3_8_port, CO => CARRYB_4_7_port, S => 
                           SUMB_4_7_port);
   S2_4_8 : FA_X1 port map( A => ab_4_8_port, B => CARRYB_3_8_port, CI => 
                           SUMB_3_9_port, CO => CARRYB_4_8_port, S => 
                           SUMB_4_8_port);
   S2_4_9 : FA_X1 port map( A => ab_4_9_port, B => CARRYB_3_9_port, CI => 
                           SUMB_3_10_port, CO => CARRYB_4_9_port, S => 
                           SUMB_4_9_port);
   S2_4_10 : FA_X1 port map( A => ab_4_10_port, B => CARRYB_3_10_port, CI => 
                           SUMB_3_11_port, CO => CARRYB_4_10_port, S => 
                           SUMB_4_10_port);
   S2_4_11 : FA_X1 port map( A => ab_4_11_port, B => CARRYB_3_11_port, CI => 
                           SUMB_3_12_port, CO => CARRYB_4_11_port, S => 
                           SUMB_4_11_port);
   S2_4_12 : FA_X1 port map( A => ab_4_12_port, B => CARRYB_3_12_port, CI => 
                           SUMB_3_13_port, CO => CARRYB_4_12_port, S => 
                           SUMB_4_12_port);
   S2_4_13 : FA_X1 port map( A => ab_4_13_port, B => CARRYB_3_13_port, CI => 
                           SUMB_3_14_port, CO => CARRYB_4_13_port, S => 
                           SUMB_4_13_port);
   S3_4_14 : FA_X1 port map( A => ab_4_14_port, B => CARRYB_3_14_port, CI => 
                           ab_3_15_port, CO => CARRYB_4_14_port, S => 
                           SUMB_4_14_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S2_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           SUMB_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S2_3_7 : FA_X1 port map( A => ab_3_7_port, B => CARRYB_2_7_port, CI => 
                           SUMB_2_8_port, CO => CARRYB_3_7_port, S => 
                           SUMB_3_7_port);
   S2_3_8 : FA_X1 port map( A => ab_3_8_port, B => CARRYB_2_8_port, CI => 
                           SUMB_2_9_port, CO => CARRYB_3_8_port, S => 
                           SUMB_3_8_port);
   S2_3_9 : FA_X1 port map( A => ab_3_9_port, B => CARRYB_2_9_port, CI => 
                           SUMB_2_10_port, CO => CARRYB_3_9_port, S => 
                           SUMB_3_9_port);
   S2_3_10 : FA_X1 port map( A => ab_3_10_port, B => CARRYB_2_10_port, CI => 
                           SUMB_2_11_port, CO => CARRYB_3_10_port, S => 
                           SUMB_3_10_port);
   S2_3_11 : FA_X1 port map( A => ab_3_11_port, B => CARRYB_2_11_port, CI => 
                           SUMB_2_12_port, CO => CARRYB_3_11_port, S => 
                           SUMB_3_11_port);
   S2_3_12 : FA_X1 port map( A => ab_3_12_port, B => CARRYB_2_12_port, CI => 
                           SUMB_2_13_port, CO => CARRYB_3_12_port, S => 
                           SUMB_3_12_port);
   S2_3_13 : FA_X1 port map( A => ab_3_13_port, B => CARRYB_2_13_port, CI => 
                           SUMB_2_14_port, CO => CARRYB_3_13_port, S => 
                           SUMB_3_13_port);
   S3_3_14 : FA_X1 port map( A => ab_3_14_port, B => CARRYB_2_14_port, CI => 
                           ab_2_15_port, CO => CARRYB_3_14_port, S => 
                           SUMB_3_14_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n30, CI => n14, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n29, CI => n9, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n26, CI => n5, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n8, CI => n28, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n25, CI => n15, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n27, CI => n13, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S2_2_6 : FA_X1 port map( A => ab_2_6_port, B => n24, CI => n12, CO => 
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   S2_2_7 : FA_X1 port map( A => ab_2_7_port, B => n23, CI => n10, CO => 
                           CARRYB_2_7_port, S => SUMB_2_7_port);
   S2_2_8 : FA_X1 port map( A => ab_2_8_port, B => n22, CI => n7, CO => 
                           CARRYB_2_8_port, S => SUMB_2_8_port);
   S2_2_9 : FA_X1 port map( A => ab_2_9_port, B => n21, CI => n11, CO => 
                           CARRYB_2_9_port, S => SUMB_2_9_port);
   S2_2_10 : FA_X1 port map( A => ab_2_10_port, B => n20, CI => n6, CO => 
                           CARRYB_2_10_port, S => SUMB_2_10_port);
   S2_2_11 : FA_X1 port map( A => ab_2_11_port, B => n19, CI => n4, CO => 
                           CARRYB_2_11_port, S => SUMB_2_11_port);
   S2_2_12 : FA_X1 port map( A => ab_2_12_port, B => n18, CI => n3, CO => 
                           CARRYB_2_12_port, S => SUMB_2_12_port);
   S2_2_13 : FA_X1 port map( A => ab_2_13_port, B => n17, CI => n2, CO => 
                           CARRYB_2_13_port, S => SUMB_2_13_port);
   S3_2_14 : FA_X1 port map( A => ab_2_14_port, B => n16, CI => ab_1_15_port, 
                           CO => CARRYB_2_14_port, S => SUMB_2_14_port);
   U2 : XOR2_X1 port map( A => ab_1_14_port, B => ab_0_15_port, Z => n2);
   U3 : XOR2_X1 port map( A => ab_1_13_port, B => ab_0_14_port, Z => n3);
   U4 : XOR2_X1 port map( A => ab_1_12_port, B => ab_0_13_port, Z => n4);
   U5 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n5);
   U6 : XOR2_X1 port map( A => ab_1_11_port, B => ab_0_12_port, Z => n6);
   U7 : XOR2_X1 port map( A => ab_1_9_port, B => ab_0_10_port, Z => n7);
   U9 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n9);
   U10 : XOR2_X1 port map( A => ab_1_8_port, B => ab_0_9_port, Z => n10);
   U11 : XOR2_X1 port map( A => ab_1_10_port, B => ab_0_11_port, Z => n11);
   U12 : XOR2_X1 port map( A => ab_1_7_port, B => ab_0_8_port, Z => n12);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n13);
   U14 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n14);
   U15 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n15);
   U28 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n28);
   U37 : XOR2_X1 port map( A => CARRYB_15_0_port, B => SUMB_15_1_port, Z => n31
                           );
   U38 : XOR2_X1 port map( A => CARRYB_15_1_port, B => SUMB_15_2_port, Z => n32
                           );
   U41 : XOR2_X1 port map( A => CARRYB_15_2_port, B => SUMB_15_3_port, Z => n35
                           );
   U43 : XOR2_X1 port map( A => CARRYB_15_3_port, B => SUMB_15_4_port, Z => n37
                           );
   U45 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U49 : XOR2_X1 port map( A => CARRYB_15_4_port, B => SUMB_15_5_port, Z => n40
                           );
   U50 : XOR2_X1 port map( A => CARRYB_15_5_port, B => SUMB_15_6_port, Z => n41
                           );
   U54 : XOR2_X1 port map( A => CARRYB_15_6_port, B => SUMB_15_7_port, Z => n43
                           );
   U56 : XOR2_X1 port map( A => CARRYB_15_7_port, B => SUMB_15_8_port, Z => n45
                           );
   U58 : XOR2_X1 port map( A => CARRYB_15_8_port, B => SUMB_15_9_port, Z => n47
                           );
   U60 : XOR2_X1 port map( A => CARRYB_15_9_port, B => SUMB_15_10_port, Z => 
                           n49);
   U62 : XOR2_X1 port map( A => CARRYB_15_10_port, B => SUMB_15_11_port, Z => 
                           n51);
   U63 : XOR2_X1 port map( A => CARRYB_15_11_port, B => SUMB_15_12_port, Z => 
                           n52);
   U67 : XOR2_X1 port map( A => CARRYB_15_12_port, B => SUMB_15_13_port, Z => 
                           n56);
   U69 : XOR2_X1 port map( A => CARRYB_15_13_port, B => SUMB_15_14_port, Z => 
                           n58);
   U71 : XOR2_X1 port map( A => CARRYB_15_14_port, B => SUMB_15_15_port, Z => 
                           n60);
   n781 <= '0';
   n782 <= '0';
   FS_1 : ALU_N32_DW01_add_1_DW01_add_3 port map( A(29) => n808, A(28) => n60, 
                           A(27) => n58, A(26) => n56, A(25) => n52, A(24) => 
                           n51, A(23) => n49, A(22) => n47, A(21) => n45, A(20)
                           => n43, A(19) => n41, A(18) => n40, A(17) => n37, 
                           A(16) => n35, A(15) => n32, A(14) => n31, A(13) => 
                           A1_13_port, A(12) => A1_12_port, A(11) => A1_11_port
                           , A(10) => A1_10_port, A(9) => A1_9_port, A(8) => 
                           A1_8_port, A(7) => A1_7_port, A(6) => A1_6_port, 
                           A(5) => A1_5_port, A(4) => A1_4_port, A(3) => 
                           A1_3_port, A(2) => A1_2_port, A(1) => A1_1_port, 
                           A(0) => A1_0_port, B(29) => n61, B(28) => n59, B(27)
                           => n57, B(26) => n55, B(25) => n54, B(24) => n53, 
                           B(23) => n50, B(22) => n48, B(21) => n46, B(20) => 
                           n44, B(19) => n42, B(18) => n38, B(17) => n36, B(16)
                           => n34, B(15) => n33, B(14) => A2_14_port, B(13) => 
                           n782, B(12) => n782, B(11) => n782, B(10) => n782, 
                           B(9) => n782, B(8) => n782, B(7) => n782, B(6) => 
                           n782, B(5) => n782, B(4) => n782, B(3) => n782, B(2)
                           => n782, B(1) => n782, B(0) => n781, CI => n781, 
                           SUM(29) => PRODUCT(31), SUM(28) => PRODUCT(30), 
                           SUM(27) => PRODUCT(29), SUM(26) => PRODUCT(28), 
                           SUM(25) => PRODUCT(27), SUM(24) => PRODUCT(26), 
                           SUM(23) => PRODUCT(25), SUM(22) => PRODUCT(24), 
                           SUM(21) => PRODUCT(23), SUM(20) => PRODUCT(22), 
                           SUM(19) => PRODUCT(21), SUM(18) => PRODUCT(20), 
                           SUM(17) => PRODUCT(19), SUM(16) => PRODUCT(18), 
                           SUM(15) => PRODUCT(17), SUM(14) => PRODUCT(16), 
                           SUM(13) => PRODUCT(15), SUM(12) => PRODUCT(14), 
                           SUM(11) => PRODUCT(13), SUM(10) => PRODUCT(12), 
                           SUM(9) => PRODUCT(11), SUM(8) => PRODUCT(10), SUM(7)
                           => PRODUCT(9), SUM(6) => PRODUCT(8), SUM(5) => 
                           PRODUCT(7), SUM(4) => PRODUCT(6), SUM(3) => 
                           PRODUCT(5), SUM(2) => PRODUCT(4), SUM(1) => 
                           PRODUCT(3), SUM(0) => PRODUCT(2), CO => n_1017);
   U17 : INV_X1 port map( A => A(1), ZN => n794);
   U18 : INV_X1 port map( A => A(0), ZN => n793);
   U19 : BUF_X1 port map( A => B(3), Z => n790);
   U20 : BUF_X1 port map( A => B(4), Z => n792);
   U21 : BUF_X1 port map( A => B(2), Z => n788);
   U22 : BUF_X1 port map( A => B(1), Z => n786);
   U23 : BUF_X1 port map( A => B(0), Z => n784);
   U24 : INV_X1 port map( A => n792, ZN => n791);
   U25 : INV_X1 port map( A => n788, ZN => n787);
   U26 : INV_X1 port map( A => n786, ZN => n785);
   U27 : INV_X1 port map( A => n790, ZN => n789);
   U29 : AND2_X1 port map( A1 => CARRYB_15_0_port, A2 => SUMB_15_1_port, ZN => 
                           n33);
   U30 : AND2_X1 port map( A1 => CARRYB_15_1_port, A2 => SUMB_15_2_port, ZN => 
                           n34);
   U31 : AND2_X1 port map( A1 => CARRYB_15_2_port, A2 => SUMB_15_3_port, ZN => 
                           n36);
   U32 : AND2_X1 port map( A1 => CARRYB_15_3_port, A2 => SUMB_15_4_port, ZN => 
                           n38);
   U33 : INV_X1 port map( A => CARRYB_15_15_port, ZN => n808);
   U34 : INV_X1 port map( A => n784, ZN => n783);
   U35 : AND2_X1 port map( A1 => CARRYB_15_14_port, A2 => SUMB_15_15_port, ZN 
                           => n61);
   U36 : NOR2_X1 port map( A1 => n819, A2 => n793, ZN => ab_0_14_port);
   U39 : NOR2_X1 port map( A1 => n818, A2 => n793, ZN => ab_0_13_port);
   U40 : NOR2_X1 port map( A1 => n817, A2 => n793, ZN => ab_0_12_port);
   U42 : NOR2_X1 port map( A1 => n816, A2 => n793, ZN => ab_0_11_port);
   U44 : NOR2_X1 port map( A1 => n815, A2 => n793, ZN => ab_0_10_port);
   U46 : NOR2_X1 port map( A1 => n814, A2 => n793, ZN => ab_0_9_port);
   U47 : NOR2_X1 port map( A1 => n813, A2 => n793, ZN => ab_0_8_port);
   U48 : NOR2_X1 port map( A1 => n812, A2 => n793, ZN => ab_0_7_port);
   U51 : NOR2_X1 port map( A1 => n811, A2 => n793, ZN => ab_0_6_port);
   U52 : NOR2_X1 port map( A1 => n810, A2 => n793, ZN => ab_0_5_port);
   U53 : NOR2_X1 port map( A1 => n791, A2 => n793, ZN => ab_0_4_port);
   U55 : NOR2_X1 port map( A1 => n789, A2 => n793, ZN => ab_0_3_port);
   U57 : NOR2_X1 port map( A1 => n787, A2 => n793, ZN => ab_0_2_port);
   U59 : NOR2_X1 port map( A1 => n785, A2 => n793, ZN => ab_0_1_port);
   U61 : NOR2_X1 port map( A1 => n819, A2 => n794, ZN => ab_1_14_port);
   U64 : NOR2_X1 port map( A1 => n818, A2 => n794, ZN => ab_1_13_port);
   U65 : NOR2_X1 port map( A1 => n817, A2 => n794, ZN => ab_1_12_port);
   U66 : NOR2_X1 port map( A1 => n816, A2 => n794, ZN => ab_1_11_port);
   U68 : NOR2_X1 port map( A1 => n815, A2 => n794, ZN => ab_1_10_port);
   U70 : NOR2_X1 port map( A1 => n814, A2 => n794, ZN => ab_1_9_port);
   U72 : NOR2_X1 port map( A1 => n813, A2 => n794, ZN => ab_1_8_port);
   U73 : NOR2_X1 port map( A1 => n812, A2 => n794, ZN => ab_1_7_port);
   U74 : NOR2_X1 port map( A1 => n811, A2 => n794, ZN => ab_1_6_port);
   U75 : NOR2_X1 port map( A1 => n810, A2 => n794, ZN => ab_1_5_port);
   U76 : NOR2_X1 port map( A1 => n791, A2 => n794, ZN => ab_1_4_port);
   U77 : NOR2_X1 port map( A1 => n789, A2 => n794, ZN => ab_1_3_port);
   U78 : NOR2_X1 port map( A1 => n787, A2 => n794, ZN => ab_1_2_port);
   U79 : NOR2_X1 port map( A1 => n785, A2 => n794, ZN => ab_1_1_port);
   U80 : NOR2_X1 port map( A1 => n783, A2 => n794, ZN => ab_1_0_port);
   U81 : NOR2_X1 port map( A1 => n783, A2 => n793, ZN => PRODUCT(0));
   U82 : NOR2_X1 port map( A1 => n786, A2 => n809, ZN => ab_15_1_port);
   U83 : NOR2_X1 port map( A1 => n784, A2 => n809, ZN => ab_15_0_port);
   U84 : NOR2_X1 port map( A1 => n790, A2 => n809, ZN => ab_15_3_port);
   U85 : NOR2_X1 port map( A1 => n788, A2 => n809, ZN => ab_15_2_port);
   U86 : NOR2_X1 port map( A1 => n792, A2 => n809, ZN => ab_15_4_port);
   U87 : AND2_X1 port map( A1 => ab_0_14_port, A2 => ab_1_13_port, ZN => n17);
   U88 : NOR2_X1 port map( A1 => n818, A2 => n795, ZN => ab_2_13_port);
   U89 : AND2_X1 port map( A1 => ab_0_13_port, A2 => ab_1_12_port, ZN => n18);
   U90 : NOR2_X1 port map( A1 => n817, A2 => n795, ZN => ab_2_12_port);
   U91 : AND2_X1 port map( A1 => ab_0_12_port, A2 => ab_1_11_port, ZN => n19);
   U92 : NOR2_X1 port map( A1 => n816, A2 => n795, ZN => ab_2_11_port);
   U93 : AND2_X1 port map( A1 => ab_0_11_port, A2 => ab_1_10_port, ZN => n20);
   U94 : NOR2_X1 port map( A1 => n815, A2 => n795, ZN => ab_2_10_port);
   U95 : AND2_X1 port map( A1 => ab_0_10_port, A2 => ab_1_9_port, ZN => n21);
   U96 : NOR2_X1 port map( A1 => n814, A2 => n795, ZN => ab_2_9_port);
   U97 : AND2_X1 port map( A1 => ab_0_9_port, A2 => ab_1_8_port, ZN => n22);
   U98 : NOR2_X1 port map( A1 => n813, A2 => n795, ZN => ab_2_8_port);
   U99 : AND2_X1 port map( A1 => ab_0_8_port, A2 => ab_1_7_port, ZN => n23);
   U100 : NOR2_X1 port map( A1 => n812, A2 => n795, ZN => ab_2_7_port);
   U101 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n24);
   U102 : NOR2_X1 port map( A1 => n811, A2 => n795, ZN => ab_2_6_port);
   U103 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n27);
   U104 : NOR2_X1 port map( A1 => n810, A2 => n795, ZN => ab_2_5_port);
   U105 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n25);
   U106 : NOR2_X1 port map( A1 => n791, A2 => n795, ZN => ab_2_4_port);
   U107 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n8);
   U108 : NOR2_X1 port map( A1 => n789, A2 => n795, ZN => ab_2_3_port);
   U109 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n26);
   U110 : NOR2_X1 port map( A1 => n787, A2 => n795, ZN => ab_2_2_port);
   U111 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n29);
   U112 : NOR2_X1 port map( A1 => n785, A2 => n795, ZN => ab_2_1_port);
   U113 : NOR2_X1 port map( A1 => n818, A2 => n796, ZN => ab_3_13_port);
   U114 : NOR2_X1 port map( A1 => n817, A2 => n796, ZN => ab_3_12_port);
   U115 : NOR2_X1 port map( A1 => n816, A2 => n796, ZN => ab_3_11_port);
   U116 : NOR2_X1 port map( A1 => n815, A2 => n796, ZN => ab_3_10_port);
   U117 : NOR2_X1 port map( A1 => n814, A2 => n796, ZN => ab_3_9_port);
   U118 : NOR2_X1 port map( A1 => n813, A2 => n796, ZN => ab_3_8_port);
   U119 : NOR2_X1 port map( A1 => n812, A2 => n796, ZN => ab_3_7_port);
   U120 : NOR2_X1 port map( A1 => n811, A2 => n796, ZN => ab_3_6_port);
   U121 : NOR2_X1 port map( A1 => n810, A2 => n796, ZN => ab_3_5_port);
   U122 : NOR2_X1 port map( A1 => n791, A2 => n796, ZN => ab_3_4_port);
   U123 : NOR2_X1 port map( A1 => n789, A2 => n796, ZN => ab_3_3_port);
   U124 : NOR2_X1 port map( A1 => n787, A2 => n796, ZN => ab_3_2_port);
   U125 : NOR2_X1 port map( A1 => n785, A2 => n796, ZN => ab_3_1_port);
   U126 : NOR2_X1 port map( A1 => n817, A2 => n797, ZN => ab_4_12_port);
   U127 : NOR2_X1 port map( A1 => n816, A2 => n797, ZN => ab_4_11_port);
   U128 : NOR2_X1 port map( A1 => n815, A2 => n797, ZN => ab_4_10_port);
   U129 : NOR2_X1 port map( A1 => n814, A2 => n797, ZN => ab_4_9_port);
   U130 : NOR2_X1 port map( A1 => n813, A2 => n797, ZN => ab_4_8_port);
   U131 : NOR2_X1 port map( A1 => n812, A2 => n797, ZN => ab_4_7_port);
   U132 : NOR2_X1 port map( A1 => n811, A2 => n797, ZN => ab_4_6_port);
   U133 : NOR2_X1 port map( A1 => n810, A2 => n797, ZN => ab_4_5_port);
   U134 : NOR2_X1 port map( A1 => n791, A2 => n797, ZN => ab_4_4_port);
   U135 : NOR2_X1 port map( A1 => n789, A2 => n797, ZN => ab_4_3_port);
   U136 : NOR2_X1 port map( A1 => n787, A2 => n797, ZN => ab_4_2_port);
   U137 : NOR2_X1 port map( A1 => n785, A2 => n797, ZN => ab_4_1_port);
   U138 : NOR2_X1 port map( A1 => n816, A2 => n798, ZN => ab_5_11_port);
   U139 : NOR2_X1 port map( A1 => n815, A2 => n798, ZN => ab_5_10_port);
   U140 : NOR2_X1 port map( A1 => n814, A2 => n798, ZN => ab_5_9_port);
   U141 : NOR2_X1 port map( A1 => n813, A2 => n798, ZN => ab_5_8_port);
   U142 : NOR2_X1 port map( A1 => n812, A2 => n798, ZN => ab_5_7_port);
   U143 : NOR2_X1 port map( A1 => n811, A2 => n798, ZN => ab_5_6_port);
   U144 : NOR2_X1 port map( A1 => n810, A2 => n798, ZN => ab_5_5_port);
   U145 : NOR2_X1 port map( A1 => n791, A2 => n798, ZN => ab_5_4_port);
   U146 : NOR2_X1 port map( A1 => n789, A2 => n798, ZN => ab_5_3_port);
   U147 : NOR2_X1 port map( A1 => n787, A2 => n798, ZN => ab_5_2_port);
   U148 : NOR2_X1 port map( A1 => n785, A2 => n798, ZN => ab_5_1_port);
   U149 : NOR2_X1 port map( A1 => n815, A2 => n799, ZN => ab_6_10_port);
   U150 : NOR2_X1 port map( A1 => n814, A2 => n799, ZN => ab_6_9_port);
   U151 : NOR2_X1 port map( A1 => n813, A2 => n799, ZN => ab_6_8_port);
   U152 : NOR2_X1 port map( A1 => n812, A2 => n799, ZN => ab_6_7_port);
   U153 : NOR2_X1 port map( A1 => n811, A2 => n799, ZN => ab_6_6_port);
   U154 : NOR2_X1 port map( A1 => n810, A2 => n799, ZN => ab_6_5_port);
   U155 : NOR2_X1 port map( A1 => n791, A2 => n799, ZN => ab_6_4_port);
   U156 : NOR2_X1 port map( A1 => n789, A2 => n799, ZN => ab_6_3_port);
   U157 : NOR2_X1 port map( A1 => n787, A2 => n799, ZN => ab_6_2_port);
   U158 : NOR2_X1 port map( A1 => n785, A2 => n799, ZN => ab_6_1_port);
   U159 : NOR2_X1 port map( A1 => n818, A2 => n797, ZN => ab_4_13_port);
   U160 : NOR2_X1 port map( A1 => n814, A2 => n800, ZN => ab_7_9_port);
   U161 : NOR2_X1 port map( A1 => n813, A2 => n800, ZN => ab_7_8_port);
   U162 : NOR2_X1 port map( A1 => n812, A2 => n800, ZN => ab_7_7_port);
   U163 : NOR2_X1 port map( A1 => n811, A2 => n800, ZN => ab_7_6_port);
   U164 : NOR2_X1 port map( A1 => n810, A2 => n800, ZN => ab_7_5_port);
   U165 : NOR2_X1 port map( A1 => n791, A2 => n800, ZN => ab_7_4_port);
   U166 : NOR2_X1 port map( A1 => n789, A2 => n800, ZN => ab_7_3_port);
   U167 : NOR2_X1 port map( A1 => n787, A2 => n800, ZN => ab_7_2_port);
   U168 : NOR2_X1 port map( A1 => n785, A2 => n800, ZN => ab_7_1_port);
   U169 : NOR2_X1 port map( A1 => n818, A2 => n798, ZN => ab_5_13_port);
   U170 : NOR2_X1 port map( A1 => n817, A2 => n798, ZN => ab_5_12_port);
   U171 : NOR2_X1 port map( A1 => n813, A2 => n801, ZN => ab_8_8_port);
   U172 : NOR2_X1 port map( A1 => n812, A2 => n801, ZN => ab_8_7_port);
   U173 : NOR2_X1 port map( A1 => n811, A2 => n801, ZN => ab_8_6_port);
   U174 : NOR2_X1 port map( A1 => n810, A2 => n801, ZN => ab_8_5_port);
   U175 : NOR2_X1 port map( A1 => n791, A2 => n801, ZN => ab_8_4_port);
   U176 : NOR2_X1 port map( A1 => n789, A2 => n801, ZN => ab_8_3_port);
   U177 : NOR2_X1 port map( A1 => n787, A2 => n801, ZN => ab_8_2_port);
   U178 : NOR2_X1 port map( A1 => n785, A2 => n801, ZN => ab_8_1_port);
   U179 : NOR2_X1 port map( A1 => n818, A2 => n799, ZN => ab_6_13_port);
   U180 : NOR2_X1 port map( A1 => n817, A2 => n799, ZN => ab_6_12_port);
   U181 : NOR2_X1 port map( A1 => n816, A2 => n799, ZN => ab_6_11_port);
   U182 : NOR2_X1 port map( A1 => n802, A2 => n812, ZN => ab_9_7_port);
   U183 : NOR2_X1 port map( A1 => n802, A2 => n811, ZN => ab_9_6_port);
   U184 : NOR2_X1 port map( A1 => n802, A2 => n810, ZN => ab_9_5_port);
   U185 : NOR2_X1 port map( A1 => n802, A2 => n791, ZN => ab_9_4_port);
   U186 : NOR2_X1 port map( A1 => n802, A2 => n789, ZN => ab_9_3_port);
   U187 : NOR2_X1 port map( A1 => n802, A2 => n787, ZN => ab_9_2_port);
   U188 : NOR2_X1 port map( A1 => n802, A2 => n785, ZN => ab_9_1_port);
   U189 : NOR2_X1 port map( A1 => n818, A2 => n800, ZN => ab_7_13_port);
   U190 : NOR2_X1 port map( A1 => n817, A2 => n800, ZN => ab_7_12_port);
   U191 : NOR2_X1 port map( A1 => n816, A2 => n800, ZN => ab_7_11_port);
   U192 : NOR2_X1 port map( A1 => n815, A2 => n800, ZN => ab_7_10_port);
   U193 : NOR2_X1 port map( A1 => n811, A2 => n803, ZN => ab_10_6_port);
   U194 : NOR2_X1 port map( A1 => n810, A2 => n803, ZN => ab_10_5_port);
   U195 : NOR2_X1 port map( A1 => n791, A2 => n803, ZN => ab_10_4_port);
   U196 : NOR2_X1 port map( A1 => n789, A2 => n803, ZN => ab_10_3_port);
   U197 : NOR2_X1 port map( A1 => n787, A2 => n803, ZN => ab_10_2_port);
   U198 : NOR2_X1 port map( A1 => n785, A2 => n803, ZN => ab_10_1_port);
   U199 : NOR2_X1 port map( A1 => n817, A2 => n801, ZN => ab_8_12_port);
   U200 : NOR2_X1 port map( A1 => n816, A2 => n801, ZN => ab_8_11_port);
   U201 : NOR2_X1 port map( A1 => n815, A2 => n801, ZN => ab_8_10_port);
   U202 : NOR2_X1 port map( A1 => n814, A2 => n801, ZN => ab_8_9_port);
   U203 : NOR2_X1 port map( A1 => n810, A2 => n804, ZN => ab_11_5_port);
   U204 : NOR2_X1 port map( A1 => n791, A2 => n804, ZN => ab_11_4_port);
   U205 : NOR2_X1 port map( A1 => n789, A2 => n804, ZN => ab_11_3_port);
   U206 : NOR2_X1 port map( A1 => n787, A2 => n804, ZN => ab_11_2_port);
   U207 : NOR2_X1 port map( A1 => n785, A2 => n804, ZN => ab_11_1_port);
   U208 : NOR2_X1 port map( A1 => n802, A2 => n816, ZN => ab_9_11_port);
   U209 : NOR2_X1 port map( A1 => n802, A2 => n815, ZN => ab_9_10_port);
   U210 : NOR2_X1 port map( A1 => n802, A2 => n814, ZN => ab_9_9_port);
   U211 : NOR2_X1 port map( A1 => n802, A2 => n813, ZN => ab_9_8_port);
   U212 : NOR2_X1 port map( A1 => n791, A2 => n805, ZN => ab_12_4_port);
   U213 : NOR2_X1 port map( A1 => n789, A2 => n805, ZN => ab_12_3_port);
   U214 : NOR2_X1 port map( A1 => n787, A2 => n805, ZN => ab_12_2_port);
   U215 : NOR2_X1 port map( A1 => n785, A2 => n805, ZN => ab_12_1_port);
   U216 : NOR2_X1 port map( A1 => n815, A2 => n803, ZN => ab_10_10_port);
   U217 : NOR2_X1 port map( A1 => n814, A2 => n803, ZN => ab_10_9_port);
   U218 : NOR2_X1 port map( A1 => n813, A2 => n803, ZN => ab_10_8_port);
   U219 : NOR2_X1 port map( A1 => n812, A2 => n803, ZN => ab_10_7_port);
   U220 : NOR2_X1 port map( A1 => n789, A2 => n806, ZN => ab_13_3_port);
   U221 : NOR2_X1 port map( A1 => n787, A2 => n806, ZN => ab_13_2_port);
   U222 : NOR2_X1 port map( A1 => n785, A2 => n806, ZN => ab_13_1_port);
   U223 : NOR2_X1 port map( A1 => n814, A2 => n804, ZN => ab_11_9_port);
   U224 : NOR2_X1 port map( A1 => n813, A2 => n804, ZN => ab_11_8_port);
   U225 : NOR2_X1 port map( A1 => n812, A2 => n804, ZN => ab_11_7_port);
   U226 : NOR2_X1 port map( A1 => n811, A2 => n804, ZN => ab_11_6_port);
   U227 : NOR2_X1 port map( A1 => n787, A2 => n807, ZN => ab_14_2_port);
   U228 : NOR2_X1 port map( A1 => n785, A2 => n807, ZN => ab_14_1_port);
   U229 : NOR2_X1 port map( A1 => n813, A2 => n805, ZN => ab_12_8_port);
   U230 : NOR2_X1 port map( A1 => n812, A2 => n805, ZN => ab_12_7_port);
   U231 : NOR2_X1 port map( A1 => n811, A2 => n805, ZN => ab_12_6_port);
   U232 : NOR2_X1 port map( A1 => n810, A2 => n805, ZN => ab_12_5_port);
   U233 : NOR2_X1 port map( A1 => n818, A2 => n801, ZN => ab_8_13_port);
   U234 : NOR2_X1 port map( A1 => n812, A2 => n806, ZN => ab_13_7_port);
   U235 : NOR2_X1 port map( A1 => n811, A2 => n806, ZN => ab_13_6_port);
   U236 : NOR2_X1 port map( A1 => n810, A2 => n806, ZN => ab_13_5_port);
   U237 : NOR2_X1 port map( A1 => n791, A2 => n806, ZN => ab_13_4_port);
   U238 : NOR2_X1 port map( A1 => n802, A2 => n818, ZN => ab_9_13_port);
   U239 : NOR2_X1 port map( A1 => n802, A2 => n817, ZN => ab_9_12_port);
   U240 : NOR2_X1 port map( A1 => n789, A2 => n807, ZN => ab_14_3_port);
   U241 : NOR2_X1 port map( A1 => n811, A2 => n807, ZN => ab_14_6_port);
   U242 : NOR2_X1 port map( A1 => n810, A2 => n807, ZN => ab_14_5_port);
   U243 : NOR2_X1 port map( A1 => n791, A2 => n807, ZN => ab_14_4_port);
   U244 : NOR2_X1 port map( A1 => n818, A2 => n803, ZN => ab_10_13_port);
   U245 : NOR2_X1 port map( A1 => n817, A2 => n803, ZN => ab_10_12_port);
   U246 : NOR2_X1 port map( A1 => n816, A2 => n803, ZN => ab_10_11_port);
   U247 : NOR2_X1 port map( A1 => n818, A2 => n804, ZN => ab_11_13_port);
   U248 : NOR2_X1 port map( A1 => n817, A2 => n804, ZN => ab_11_12_port);
   U249 : NOR2_X1 port map( A1 => n816, A2 => n804, ZN => ab_11_11_port);
   U250 : NOR2_X1 port map( A1 => n815, A2 => n804, ZN => ab_11_10_port);
   U251 : NOR2_X1 port map( A1 => n817, A2 => n805, ZN => ab_12_12_port);
   U252 : NOR2_X1 port map( A1 => n816, A2 => n805, ZN => ab_12_11_port);
   U253 : NOR2_X1 port map( A1 => n815, A2 => n805, ZN => ab_12_10_port);
   U254 : NOR2_X1 port map( A1 => n814, A2 => n805, ZN => ab_12_9_port);
   U255 : NOR2_X1 port map( A1 => n816, A2 => n806, ZN => ab_13_11_port);
   U256 : NOR2_X1 port map( A1 => n815, A2 => n806, ZN => ab_13_10_port);
   U257 : NOR2_X1 port map( A1 => n814, A2 => n806, ZN => ab_13_9_port);
   U258 : NOR2_X1 port map( A1 => n813, A2 => n806, ZN => ab_13_8_port);
   U259 : NOR2_X1 port map( A1 => n812, A2 => n807, ZN => ab_14_7_port);
   U260 : NOR2_X1 port map( A1 => n815, A2 => n807, ZN => ab_14_10_port);
   U261 : NOR2_X1 port map( A1 => n814, A2 => n807, ZN => ab_14_9_port);
   U262 : NOR2_X1 port map( A1 => n813, A2 => n807, ZN => ab_14_8_port);
   U263 : NOR2_X1 port map( A1 => n818, A2 => n805, ZN => ab_12_13_port);
   U264 : NOR2_X1 port map( A1 => n817, A2 => n806, ZN => ab_13_12_port);
   U265 : NOR2_X1 port map( A1 => n816, A2 => n807, ZN => ab_14_11_port);
   U266 : NOR2_X1 port map( A1 => n818, A2 => n806, ZN => ab_13_13_port);
   U267 : NOR2_X1 port map( A1 => n817, A2 => n807, ZN => ab_14_12_port);
   U268 : NOR2_X1 port map( A1 => n818, A2 => n807, ZN => ab_14_13_port);
   U269 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n30);
   U270 : NOR2_X1 port map( A1 => n783, A2 => n795, ZN => ab_2_0_port);
   U271 : NOR2_X1 port map( A1 => n783, A2 => n796, ZN => ab_3_0_port);
   U272 : NOR2_X1 port map( A1 => n783, A2 => n797, ZN => ab_4_0_port);
   U273 : NOR2_X1 port map( A1 => n783, A2 => n798, ZN => ab_5_0_port);
   U274 : NOR2_X1 port map( A1 => n783, A2 => n799, ZN => ab_6_0_port);
   U275 : NOR2_X1 port map( A1 => n783, A2 => n800, ZN => ab_7_0_port);
   U276 : NOR2_X1 port map( A1 => n783, A2 => n801, ZN => ab_8_0_port);
   U277 : NOR2_X1 port map( A1 => n802, A2 => n783, ZN => ab_9_0_port);
   U278 : NOR2_X1 port map( A1 => n783, A2 => n803, ZN => ab_10_0_port);
   U279 : NOR2_X1 port map( A1 => n783, A2 => n804, ZN => ab_11_0_port);
   U280 : NOR2_X1 port map( A1 => n783, A2 => n805, ZN => ab_12_0_port);
   U281 : NOR2_X1 port map( A1 => n783, A2 => n806, ZN => ab_13_0_port);
   U282 : NOR2_X1 port map( A1 => n783, A2 => n807, ZN => ab_14_0_port);
   U283 : NOR2_X1 port map( A1 => n820, A2 => n809, ZN => ab_15_15_port);
   U284 : AND2_X1 port map( A1 => CARRYB_15_4_port, A2 => SUMB_15_5_port, ZN =>
                           n42);
   U285 : AND2_X1 port map( A1 => CARRYB_15_5_port, A2 => SUMB_15_6_port, ZN =>
                           n44);
   U286 : AND2_X1 port map( A1 => CARRYB_15_6_port, A2 => SUMB_15_7_port, ZN =>
                           n46);
   U287 : AND2_X1 port map( A1 => CARRYB_15_8_port, A2 => SUMB_15_9_port, ZN =>
                           n50);
   U288 : AND2_X1 port map( A1 => CARRYB_15_9_port, A2 => SUMB_15_10_port, ZN 
                           => n53);
   U289 : AND2_X1 port map( A1 => CARRYB_15_10_port, A2 => SUMB_15_11_port, ZN 
                           => n54);
   U290 : AND2_X1 port map( A1 => CARRYB_15_12_port, A2 => SUMB_15_13_port, ZN 
                           => n57);
   U291 : AND2_X1 port map( A1 => CARRYB_15_13_port, A2 => SUMB_15_14_port, ZN 
                           => n59);
   U292 : AND2_X1 port map( A1 => CARRYB_15_7_port, A2 => SUMB_15_8_port, ZN =>
                           n48);
   U293 : AND2_X1 port map( A1 => CARRYB_15_11_port, A2 => SUMB_15_12_port, ZN 
                           => n55);
   U294 : INV_X1 port map( A => A(15), ZN => n809);
   U295 : INV_X1 port map( A => A(3), ZN => n796);
   U296 : INV_X1 port map( A => A(4), ZN => n797);
   U297 : INV_X1 port map( A => A(5), ZN => n798);
   U298 : INV_X1 port map( A => A(6), ZN => n799);
   U299 : INV_X1 port map( A => A(7), ZN => n800);
   U300 : INV_X1 port map( A => A(8), ZN => n801);
   U301 : INV_X1 port map( A => A(10), ZN => n803);
   U302 : INV_X1 port map( A => A(11), ZN => n804);
   U303 : INV_X1 port map( A => A(12), ZN => n805);
   U304 : INV_X1 port map( A => A(13), ZN => n806);
   U305 : INV_X1 port map( A => A(14), ZN => n807);
   U306 : INV_X1 port map( A => A(2), ZN => n795);
   U307 : INV_X1 port map( A => A(9), ZN => n802);
   U308 : INV_X1 port map( A => B(15), ZN => n820);
   U309 : INV_X1 port map( A => B(14), ZN => n819);
   U310 : INV_X1 port map( A => B(13), ZN => n818);
   U311 : INV_X1 port map( A => B(12), ZN => n817);
   U312 : INV_X1 port map( A => B(11), ZN => n816);
   U313 : INV_X1 port map( A => B(10), ZN => n815);
   U314 : INV_X1 port map( A => B(9), ZN => n814);
   U315 : INV_X1 port map( A => B(8), ZN => n813);
   U316 : INV_X1 port map( A => B(7), ZN => n812);
   U317 : INV_X1 port map( A => B(6), ZN => n811);
   U318 : INV_X1 port map( A => B(5), ZN => n810);
   U319 : NOR2_X1 port map( A1 => A(0), A2 => n820, ZN => ab_0_15_port);
   U320 : NOR2_X1 port map( A1 => B(5), A2 => n809, ZN => ab_15_5_port);
   U321 : NOR2_X1 port map( A1 => B(7), A2 => n809, ZN => ab_15_7_port);
   U322 : NOR2_X1 port map( A1 => B(6), A2 => n809, ZN => ab_15_6_port);
   U323 : NOR2_X1 port map( A1 => B(9), A2 => n809, ZN => ab_15_9_port);
   U324 : NOR2_X1 port map( A1 => B(8), A2 => n809, ZN => ab_15_8_port);
   U325 : NOR2_X1 port map( A1 => B(10), A2 => n809, ZN => ab_15_10_port);
   U326 : NOR2_X1 port map( A1 => B(11), A2 => n809, ZN => ab_15_11_port);
   U327 : NOR2_X1 port map( A1 => B(12), A2 => n809, ZN => ab_15_12_port);
   U328 : NOR2_X1 port map( A1 => B(13), A2 => n809, ZN => ab_15_13_port);
   U329 : NOR2_X1 port map( A1 => A(14), A2 => n820, ZN => ab_14_15_port);
   U330 : NOR2_X1 port map( A1 => B(14), A2 => n809, ZN => ab_15_14_port);
   U331 : AND2_X1 port map( A1 => ab_0_15_port, A2 => ab_1_14_port, ZN => n16);
   U332 : NOR2_X1 port map( A1 => A(1), A2 => n820, ZN => ab_1_15_port);
   U333 : NOR2_X1 port map( A1 => n819, A2 => n795, ZN => ab_2_14_port);
   U334 : NOR2_X1 port map( A1 => A(2), A2 => n820, ZN => ab_2_15_port);
   U335 : NOR2_X1 port map( A1 => n819, A2 => n796, ZN => ab_3_14_port);
   U336 : NOR2_X1 port map( A1 => A(3), A2 => n820, ZN => ab_3_15_port);
   U337 : NOR2_X1 port map( A1 => n819, A2 => n797, ZN => ab_4_14_port);
   U338 : NOR2_X1 port map( A1 => A(4), A2 => n820, ZN => ab_4_15_port);
   U339 : NOR2_X1 port map( A1 => n819, A2 => n798, ZN => ab_5_14_port);
   U340 : NOR2_X1 port map( A1 => A(5), A2 => n820, ZN => ab_5_15_port);
   U341 : NOR2_X1 port map( A1 => n819, A2 => n799, ZN => ab_6_14_port);
   U342 : NOR2_X1 port map( A1 => A(6), A2 => n820, ZN => ab_6_15_port);
   U343 : NOR2_X1 port map( A1 => n819, A2 => n800, ZN => ab_7_14_port);
   U344 : NOR2_X1 port map( A1 => A(7), A2 => n820, ZN => ab_7_15_port);
   U345 : NOR2_X1 port map( A1 => n819, A2 => n801, ZN => ab_8_14_port);
   U346 : NOR2_X1 port map( A1 => A(8), A2 => n820, ZN => ab_8_15_port);
   U347 : NOR2_X1 port map( A1 => n802, A2 => n819, ZN => ab_9_14_port);
   U348 : NOR2_X1 port map( A1 => A(9), A2 => n820, ZN => ab_9_15_port);
   U349 : NOR2_X1 port map( A1 => n819, A2 => n803, ZN => ab_10_14_port);
   U350 : NOR2_X1 port map( A1 => A(10), A2 => n820, ZN => ab_10_15_port);
   U351 : NOR2_X1 port map( A1 => n819, A2 => n804, ZN => ab_11_14_port);
   U352 : NOR2_X1 port map( A1 => A(11), A2 => n820, ZN => ab_11_15_port);
   U353 : NOR2_X1 port map( A1 => n819, A2 => n805, ZN => ab_12_14_port);
   U354 : NOR2_X1 port map( A1 => A(12), A2 => n820, ZN => ab_12_15_port);
   U355 : NOR2_X1 port map( A1 => n819, A2 => n806, ZN => ab_13_14_port);
   U356 : NOR2_X1 port map( A1 => A(13), A2 => n820, ZN => ab_13_15_port);
   U357 : NOR2_X1 port map( A1 => n819, A2 => n807, ZN => ab_14_14_port);

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_N32_DW01_sub_0;

architecture SYN_rpl of ALU_N32_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n580, n581, n582,
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n_1020 : std_logic;

begin
   
   U2_31 : FA_X1 port map( A => A(31), B => n611, CI => carry_31_port, CO => 
                           n_1020, S => DIFF(31));
   U2_30 : FA_X1 port map( A => A(30), B => n610, CI => carry_30_port, CO => 
                           carry_31_port, S => DIFF(30));
   U2_29 : FA_X1 port map( A => A(29), B => n609, CI => carry_29_port, CO => 
                           carry_30_port, S => DIFF(29));
   U2_28 : FA_X1 port map( A => A(28), B => n608, CI => carry_28_port, CO => 
                           carry_29_port, S => DIFF(28));
   U2_27 : FA_X1 port map( A => A(27), B => n607, CI => carry_27_port, CO => 
                           carry_28_port, S => DIFF(27));
   U2_26 : FA_X1 port map( A => A(26), B => n606, CI => carry_26_port, CO => 
                           carry_27_port, S => DIFF(26));
   U2_25 : FA_X1 port map( A => A(25), B => n605, CI => carry_25_port, CO => 
                           carry_26_port, S => DIFF(25));
   U2_24 : FA_X1 port map( A => A(24), B => n604, CI => carry_24_port, CO => 
                           carry_25_port, S => DIFF(24));
   U2_23 : FA_X1 port map( A => A(23), B => n603, CI => carry_23_port, CO => 
                           carry_24_port, S => DIFF(23));
   U2_22 : FA_X1 port map( A => A(22), B => n602, CI => carry_22_port, CO => 
                           carry_23_port, S => DIFF(22));
   U2_21 : FA_X1 port map( A => A(21), B => n601, CI => carry_21_port, CO => 
                           carry_22_port, S => DIFF(21));
   U2_20 : FA_X1 port map( A => A(20), B => n600, CI => carry_20_port, CO => 
                           carry_21_port, S => DIFF(20));
   U2_19 : FA_X1 port map( A => A(19), B => n599, CI => carry_19_port, CO => 
                           carry_20_port, S => DIFF(19));
   U2_18 : FA_X1 port map( A => A(18), B => n598, CI => carry_18_port, CO => 
                           carry_19_port, S => DIFF(18));
   U2_17 : FA_X1 port map( A => A(17), B => n597, CI => carry_17_port, CO => 
                           carry_18_port, S => DIFF(17));
   U2_16 : FA_X1 port map( A => A(16), B => n596, CI => carry_16_port, CO => 
                           carry_17_port, S => DIFF(16));
   U2_15 : FA_X1 port map( A => A(15), B => n595, CI => carry_15_port, CO => 
                           carry_16_port, S => DIFF(15));
   U2_14 : FA_X1 port map( A => A(14), B => n594, CI => carry_14_port, CO => 
                           carry_15_port, S => DIFF(14));
   U2_13 : FA_X1 port map( A => A(13), B => n593, CI => carry_13_port, CO => 
                           carry_14_port, S => DIFF(13));
   U2_12 : FA_X1 port map( A => A(12), B => n592, CI => carry_12_port, CO => 
                           carry_13_port, S => DIFF(12));
   U2_11 : FA_X1 port map( A => A(11), B => n591, CI => carry_11_port, CO => 
                           carry_12_port, S => DIFF(11));
   U2_10 : FA_X1 port map( A => A(10), B => n590, CI => carry_10_port, CO => 
                           carry_11_port, S => DIFF(10));
   U2_9 : FA_X1 port map( A => A(9), B => n589, CI => carry_9_port, CO => 
                           carry_10_port, S => DIFF(9));
   U2_8 : FA_X1 port map( A => A(8), B => n588, CI => carry_8_port, CO => 
                           carry_9_port, S => DIFF(8));
   U2_7 : FA_X1 port map( A => A(7), B => n587, CI => carry_7_port, CO => 
                           carry_8_port, S => DIFF(7));
   U2_6 : FA_X1 port map( A => A(6), B => n586, CI => carry_6_port, CO => 
                           carry_7_port, S => DIFF(6));
   U2_5 : FA_X1 port map( A => A(5), B => n585, CI => carry_5_port, CO => 
                           carry_6_port, S => DIFF(5));
   U2_4 : FA_X1 port map( A => A(4), B => n583, CI => carry_4_port, CO => 
                           carry_5_port, S => DIFF(4));
   U2_3 : FA_X1 port map( A => A(3), B => n582, CI => carry_3_port, CO => 
                           carry_4_port, S => DIFF(3));
   U2_2 : FA_X1 port map( A => A(2), B => n581, CI => carry_2_port, CO => 
                           carry_3_port, S => DIFF(2));
   U2_1 : FA_X1 port map( A => A(1), B => n580, CI => carry_1_port, CO => 
                           carry_2_port, S => DIFF(1));
   U33 : XOR2_X1 port map( A => B(0), B => A(0), Z => DIFF(0));
   U1 : INV_X1 port map( A => B(1), ZN => n580);
   U2 : NAND2_X1 port map( A1 => B(0), A2 => n584, ZN => carry_1_port);
   U3 : INV_X1 port map( A => A(0), ZN => n584);
   U4 : INV_X1 port map( A => B(2), ZN => n581);
   U5 : INV_X1 port map( A => B(3), ZN => n582);
   U6 : INV_X1 port map( A => B(4), ZN => n583);
   U7 : INV_X1 port map( A => B(5), ZN => n585);
   U8 : INV_X1 port map( A => B(6), ZN => n586);
   U9 : INV_X1 port map( A => B(7), ZN => n587);
   U10 : INV_X1 port map( A => B(8), ZN => n588);
   U11 : INV_X1 port map( A => B(9), ZN => n589);
   U12 : INV_X1 port map( A => B(10), ZN => n590);
   U13 : INV_X1 port map( A => B(11), ZN => n591);
   U14 : INV_X1 port map( A => B(12), ZN => n592);
   U15 : INV_X1 port map( A => B(13), ZN => n593);
   U16 : INV_X1 port map( A => B(14), ZN => n594);
   U17 : INV_X1 port map( A => B(15), ZN => n595);
   U18 : INV_X1 port map( A => B(16), ZN => n596);
   U19 : INV_X1 port map( A => B(17), ZN => n597);
   U20 : INV_X1 port map( A => B(18), ZN => n598);
   U21 : INV_X1 port map( A => B(19), ZN => n599);
   U22 : INV_X1 port map( A => B(20), ZN => n600);
   U23 : INV_X1 port map( A => B(21), ZN => n601);
   U24 : INV_X1 port map( A => B(22), ZN => n602);
   U25 : INV_X1 port map( A => B(23), ZN => n603);
   U26 : INV_X1 port map( A => B(24), ZN => n604);
   U27 : INV_X1 port map( A => B(25), ZN => n605);
   U28 : INV_X1 port map( A => B(26), ZN => n606);
   U29 : INV_X1 port map( A => B(27), ZN => n607);
   U30 : INV_X1 port map( A => B(28), ZN => n608);
   U31 : INV_X1 port map( A => B(29), ZN => n609);
   U32 : INV_X1 port map( A => B(30), ZN => n610);
   U34 : INV_X1 port map( A => B(31), ZN => n611);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_N32_DW01_add_0;

architecture SYN_rpl of ALU_N32_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1023 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1023, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end ALU_N32_DW01_ash_0;

architecture SYN_mx2 of ALU_N32_DW01_ash_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, n24, n25, n26, n27, n28, n29, n30, n31, n462, n463, n464
      , n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487 : 
      std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n478, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n478, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n478, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n478, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n478, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n478, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => SH(4), Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => SH(4), Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => n487, S => SH(4), Z 
                           => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => n483, S => SH(4), Z 
                           => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => n485, S => SH(4), Z 
                           => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => n481, S => n478, Z 
                           => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => n486, S => SH(4), Z 
                           => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n482, S => SH(4), Z 
                           => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => n484, S => SH(4), Z 
                           => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => n480, S => SH(4), Z 
                           => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n474, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => SH(3), Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => SH(3), Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n474, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n474, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n474, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n474, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n474, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n474, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n474, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n474, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n474, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n474, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n474, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n474, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n474, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n474, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n474, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n474, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           SH(3), Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n470, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n470, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n470, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n470, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n470, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n470, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n470, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n470, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n470, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n470, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n470, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n470, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n470, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n470, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n470, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n470, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n470, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n466, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n466, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n466, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n466, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n466, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n466, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n466, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n466, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n466, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n466, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n466, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n466, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n466, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n466, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n466, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n466, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n466, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n466, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n463, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n463, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n463, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n462, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n463, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n462, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n463, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n462, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n463, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n463, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n463, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n463, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n463, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n463, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n463, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n462, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n463, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n462, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n462, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n462, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n462, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n462, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n462, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n462, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n462, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n462, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n462, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n463, Z => 
                           ML_int_1_1_port);
   U3 : BUF_X1 port map( A => n469, Z => n467);
   U4 : BUF_X1 port map( A => n473, Z => n471);
   U5 : BUF_X1 port map( A => n477, Z => n475);
   U6 : BUF_X1 port map( A => n465, Z => n464);
   U7 : NOR2_X1 port map( A1 => n478, A2 => n31, ZN => B(0));
   U8 : INV_X1 port map( A => n467, ZN => n466);
   U9 : INV_X1 port map( A => n471, ZN => n470);
   U10 : INV_X1 port map( A => n475, ZN => n474);
   U11 : INV_X1 port map( A => n27, ZN => n481);
   U12 : INV_X1 port map( A => n26, ZN => n485);
   U13 : INV_X1 port map( A => n25, ZN => n483);
   U14 : INV_X1 port map( A => n24, ZN => n487);
   U15 : INV_X1 port map( A => n31, ZN => n480);
   U16 : INV_X1 port map( A => n30, ZN => n484);
   U17 : INV_X1 port map( A => n29, ZN => n482);
   U18 : INV_X1 port map( A => n28, ZN => n486);
   U19 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n476, ZN => n31);
   U20 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n476, ZN => n30);
   U21 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n476, ZN => n29);
   U22 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n476, ZN => n28);
   U23 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n476, ZN => n27);
   U24 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n476, ZN => n26);
   U25 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n476, ZN => n25);
   U26 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n476, ZN => n24);
   U27 : INV_X1 port map( A => n479, ZN => n478);
   U28 : BUF_X1 port map( A => n477, Z => n476);
   U29 : INV_X1 port map( A => n464, ZN => n462);
   U30 : INV_X1 port map( A => n464, ZN => n463);
   U31 : BUF_X1 port map( A => n473, Z => n472);
   U32 : BUF_X1 port map( A => n469, Z => n468);
   U33 : INV_X1 port map( A => SH(4), ZN => n479);
   U34 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n472, ZN => 
                           ML_int_3_2_port);
   U35 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n472, ZN => 
                           ML_int_3_3_port);
   U36 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n472, ZN => 
                           ML_int_3_0_port);
   U37 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n472, ZN => 
                           ML_int_3_1_port);
   U38 : INV_X1 port map( A => SH(1), ZN => n469);
   U39 : INV_X1 port map( A => SH(2), ZN => n473);
   U40 : INV_X1 port map( A => SH(3), ZN => n477);
   U41 : NOR2_X1 port map( A1 => n478, A2 => n30, ZN => B(1));
   U42 : NOR2_X1 port map( A1 => n478, A2 => n29, ZN => B(2));
   U43 : NOR2_X1 port map( A1 => n478, A2 => n28, ZN => B(3));
   U44 : NOR2_X1 port map( A1 => n478, A2 => n27, ZN => B(4));
   U45 : NOR2_X1 port map( A1 => n478, A2 => n26, ZN => B(5));
   U46 : NOR2_X1 port map( A1 => n478, A2 => n25, ZN => B(6));
   U47 : NOR2_X1 port map( A1 => n478, A2 => n24, ZN => B(7));
   U48 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n479, ZN => B(8));
   U49 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n479, ZN => B(9));
   U50 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n479, ZN => B(10));
   U51 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n479, ZN => B(11));
   U52 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n479, ZN => B(12));
   U53 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n479, ZN => B(13));
   U54 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n479, ZN => B(14));
   U55 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n479, ZN => B(15));
   U56 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n468, ZN => 
                           ML_int_2_1_port);
   U57 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n468, ZN => 
                           ML_int_2_0_port);
   U58 : INV_X1 port map( A => SH(0), ZN => n465);
   U59 : AND2_X1 port map( A1 => A(0), A2 => n465, ZN => ML_int_1_0_port);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end ALU_N32_DW_sra_0;

architecture SYN_mx2 of ALU_N32_DW_sra_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n1198, n1199,
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : NOR2_X2 port map( A1 => n1201, A2 => SH(3), ZN => n112);
   U28 : NOR2_X2 port map( A1 => n1198, A2 => n1199, ZN => n95);
   U177 : MUX2_X1 port map( A => A(30), B => A(31), S => n98, Z => n123);
   U3 : NOR2_X2 port map( A1 => n1200, A2 => SH(3), ZN => n114);
   U4 : NAND2_X1 port map( A1 => n1205, A2 => A(31), ZN => n100);
   U5 : BUF_X1 port map( A => n1202, Z => n1204);
   U6 : INV_X1 port map( A => n97, ZN => n1254);
   U7 : INV_X1 port map( A => n94, ZN => n1255);
   U8 : INV_X1 port map( A => n88, ZN => n1256);
   U9 : INV_X1 port map( A => n61, ZN => n1257);
   U10 : INV_X1 port map( A => n1204, ZN => n1203);
   U11 : INV_X1 port map( A => n98, ZN => n1253);
   U12 : NOR2_X2 port map( A1 => n1199, A2 => SH(0), ZN => n94);
   U13 : NAND2_X1 port map( A1 => n114, A2 => n1203, ZN => n61);
   U14 : AND2_X1 port map( A1 => n1200, A2 => n166, ZN => n66);
   U15 : INV_X1 port map( A => n95, ZN => n1252);
   U16 : NAND2_X1 port map( A1 => SH(0), A2 => n1199, ZN => n97);
   U17 : NAND2_X1 port map( A1 => n112, A2 => n1203, ZN => n88);
   U18 : AND2_X1 port map( A1 => n166, A2 => n1201, ZN => n64);
   U19 : BUF_X1 port map( A => n1202, Z => n1205);
   U20 : INV_X1 port map( A => n1200, ZN => n1201);
   U21 : NAND2_X1 port map( A1 => n1198, A2 => n1199, ZN => n98);
   U22 : AND2_X1 port map( A1 => SH(3), A2 => n1201, ZN => n122);
   U23 : AOI21_X1 port map( B1 => n111, B2 => n114, A => n143, ZN => n107);
   U24 : AND2_X1 port map( A1 => n1200, A2 => SH(3), ZN => n136);
   U25 : AND2_X1 port map( A1 => SH(3), A2 => n1203, ZN => n166);
   U26 : BUF_X1 port map( A => SH(2), Z => n1200);
   U27 : BUF_X1 port map( A => SH(4), Z => n1202);
   U29 : INV_X1 port map( A => SH(1), ZN => n1199);
   U30 : OAI222_X1 port map( A1 => n98, A2 => n1246, B1 => n97, B2 => n1247, C1
                           => n1199, C2 => n1249, ZN => n111);
   U31 : AOI221_X1 port map( B1 => n72, B2 => n112, C1 => n71, C2 => n114, A =>
                           n1237, ZN => n139);
   U32 : INV_X1 port map( A => n169, ZN => n1237);
   U33 : AOI22_X1 port map( A1 => n136, A2 => n115, B1 => n122, B2 => n116, ZN 
                           => n169);
   U34 : AOI221_X1 port map( B1 => n67, B2 => n112, C1 => n65, C2 => n114, A =>
                           n1239, ZN => n127);
   U35 : INV_X1 port map( A => n138, ZN => n1239);
   U36 : AOI22_X1 port map( A1 => n136, A2 => n111, B1 => n122, B2 => n113, ZN 
                           => n138);
   U37 : AOI221_X1 port map( B1 => n123, B2 => n136, C1 => n119, C2 => n122, A 
                           => n1229, ZN => n101);
   U38 : INV_X1 port map( A => n137, ZN => n1229);
   U39 : AOI22_X1 port map( A1 => n112, A2 => n120, B1 => n114, B2 => n81, ZN 
                           => n137);
   U40 : AOI221_X1 port map( B1 => n118, B2 => n112, C1 => n77, C2 => n114, A 
                           => n1242, ZN => n89);
   U41 : INV_X1 port map( A => n134, ZN => n1242);
   U42 : AOI21_X1 port map( B1 => n122, B2 => n117, A => n124, ZN => n134);
   U43 : AOI221_X1 port map( B1 => n116, B2 => n112, C1 => n72, C2 => n114, A 
                           => n1244, ZN => n86);
   U44 : INV_X1 port map( A => n126, ZN => n1244);
   U45 : AOI21_X1 port map( B1 => n122, B2 => n115, A => n124, ZN => n126);
   U46 : AOI221_X1 port map( B1 => n113, B2 => n112, C1 => n67, C2 => n114, A 
                           => n1245, ZN => n83);
   U47 : INV_X1 port map( A => n125, ZN => n1245);
   U48 : AOI21_X1 port map( B1 => n122, B2 => n111, A => n124, ZN => n125);
   U49 : AOI221_X1 port map( B1 => n119, B2 => n112, C1 => n120, C2 => n114, A 
                           => n1248, ZN => n79);
   U50 : INV_X1 port map( A => n121, ZN => n1248);
   U51 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n121);
   U52 : AOI221_X1 port map( B1 => n117, B2 => n112, C1 => n118, C2 => n114, A 
                           => n1251, ZN => n74);
   U53 : AOI221_X1 port map( B1 => n115, B2 => n112, C1 => n116, C2 => n114, A 
                           => n1251, ZN => n69);
   U54 : AOI221_X1 port map( B1 => n111, B2 => n112, C1 => n113, C2 => n114, A 
                           => n1251, ZN => n62);
   U55 : AOI221_X1 port map( B1 => n123, B2 => n112, C1 => n119, C2 => n114, A 
                           => n1251, ZN => n110);
   U56 : OAI21_X1 port map( B1 => n1201, B2 => n1249, A => n135, ZN => n143);
   U57 : NOR2_X1 port map( A1 => n135, A2 => n1201, ZN => n124);
   U58 : OAI221_X1 port map( B1 => n85, B2 => n61, C1 => n86, C2 => n1203, A =>
                           n87, ZN => B_4_port);
   U59 : AOI222_X1 port map( A1 => n1256, A2 => n1212, B1 => n64, B2 => n1221, 
                           C1 => n66, C2 => n71, ZN => n87);
   U60 : OAI221_X1 port map( B1 => n82, B2 => n61, C1 => n83, C2 => n1203, A =>
                           n84, ZN => B_5_port);
   U61 : AOI222_X1 port map( A1 => n1256, A2 => n1214, B1 => n64, B2 => n1223, 
                           C1 => n66, C2 => n65, ZN => n84);
   U62 : OAI221_X1 port map( B1 => n78, B2 => n61, C1 => n79, C2 => n1203, A =>
                           n80, ZN => B_6_port);
   U63 : AOI222_X1 port map( A1 => n1256, A2 => n1216, B1 => n64, B2 => n1225, 
                           C1 => n66, C2 => n81, ZN => n80);
   U64 : OAI221_X1 port map( B1 => n73, B2 => n61, C1 => n74, C2 => n1203, A =>
                           n75, ZN => B_7_port);
   U65 : AOI222_X1 port map( A1 => n1256, A2 => n1218, B1 => n64, B2 => n76, C1
                           => n66, C2 => n77, ZN => n75);
   U66 : OAI221_X1 port map( B1 => n68, B2 => n61, C1 => n69, C2 => n1203, A =>
                           n70, ZN => B_8_port);
   U67 : AOI222_X1 port map( A1 => n1256, A2 => n1221, B1 => n64, B2 => n71, C1
                           => n66, C2 => n72, ZN => n70);
   U68 : OAI221_X1 port map( B1 => n60, B2 => n61, C1 => n62, C2 => n1203, A =>
                           n63, ZN => B_9_port);
   U69 : AOI222_X1 port map( A1 => n1256, A2 => n1223, B1 => n64, B2 => n65, C1
                           => n66, C2 => n67, ZN => n63);
   U70 : OAI221_X1 port map( B1 => n104, B2 => n61, C1 => n110, C2 => n1203, A 
                           => n157, ZN => B_10_port);
   U71 : AOI222_X1 port map( A1 => n1256, A2 => n1225, B1 => n64, B2 => n81, C1
                           => n66, C2 => n120, ZN => n157);
   U72 : OAI221_X1 port map( B1 => n92, B2 => n61, C1 => n109, C2 => n1203, A 
                           => n151, ZN => B_11_port);
   U73 : AOI222_X1 port map( A1 => n1256, A2 => n76, B1 => n64, B2 => n77, C1 
                           => n66, C2 => n118, ZN => n151);
   U74 : OAI221_X1 port map( B1 => n149, B2 => n61, C1 => n108, C2 => n1203, A 
                           => n150, ZN => B_12_port);
   U75 : AOI222_X1 port map( A1 => n1256, A2 => n71, B1 => n64, B2 => n72, C1 
                           => n66, C2 => n116, ZN => n150);
   U76 : OAI221_X1 port map( B1 => n132, B2 => n61, C1 => n107, C2 => n1203, A 
                           => n144, ZN => B_13_port);
   U77 : AOI222_X1 port map( A1 => n1256, A2 => n65, B1 => n64, B2 => n67, C1 
                           => n66, C2 => n113, ZN => n144);
   U78 : OAI221_X1 port map( B1 => n141, B2 => n61, C1 => n99, C2 => n1203, A 
                           => n142, ZN => B_14_port);
   U79 : AOI222_X1 port map( A1 => n1256, A2 => n81, B1 => n64, B2 => n120, C1 
                           => n66, C2 => n119, ZN => n142);
   U80 : OAI221_X1 port map( B1 => n1231, B2 => n88, C1 => n1227, C2 => n61, A 
                           => n140, ZN => B_15_port);
   U81 : INV_X1 port map( A => n76, ZN => n1227);
   U82 : INV_X1 port map( A => n77, ZN => n1231);
   U83 : AOI221_X1 port map( B1 => n66, B2 => n117, C1 => n64, C2 => n118, A =>
                           n1250, ZN => n140);
   U84 : AOI21_X1 port map( B1 => n117, B2 => n114, A => n143, ZN => n109);
   U85 : AOI21_X1 port map( B1 => n115, B2 => n114, A => n143, ZN => n108);
   U86 : AOI21_X1 port map( B1 => n123, B2 => n114, A => n143, ZN => n99);
   U87 : OAI21_X1 port map( B1 => n1205, B2 => n139, A => n100, ZN => B_16_port
                           );
   U88 : OAI21_X1 port map( B1 => n1205, B2 => n127, A => n100, ZN => B_17_port
                           );
   U89 : OAI21_X1 port map( B1 => n1204, B2 => n101, A => n100, ZN => B_18_port
                           );
   U90 : OAI21_X1 port map( B1 => n1204, B2 => n89, A => n100, ZN => B_19_port)
                           ;
   U91 : OAI21_X1 port map( B1 => n1204, B2 => n86, A => n100, ZN => B_20_port)
                           ;
   U92 : OAI21_X1 port map( B1 => n1204, B2 => n83, A => n100, ZN => B_21_port)
                           ;
   U93 : OAI21_X1 port map( B1 => n1204, B2 => n79, A => n100, ZN => B_22_port)
                           ;
   U94 : OAI21_X1 port map( B1 => n1204, B2 => n74, A => n100, ZN => B_23_port)
                           ;
   U95 : OAI21_X1 port map( B1 => n1204, B2 => n69, A => n100, ZN => B_24_port)
                           ;
   U96 : OAI21_X1 port map( B1 => n1204, B2 => n62, A => n100, ZN => B_25_port)
                           ;
   U97 : OAI21_X1 port map( B1 => n1204, B2 => n110, A => n100, ZN => B_26_port
                           );
   U98 : OAI21_X1 port map( B1 => n1204, B2 => n109, A => n100, ZN => B_27_port
                           );
   U99 : OAI21_X1 port map( B1 => n1204, B2 => n108, A => n100, ZN => B_28_port
                           );
   U100 : OAI21_X1 port map( B1 => n1204, B2 => n107, A => n100, ZN => 
                           B_29_port);
   U101 : OAI21_X1 port map( B1 => n1204, B2 => n99, A => n100, ZN => B_30_port
                           );
   U102 : INV_X1 port map( A => n149, ZN => n1221);
   U103 : INV_X1 port map( A => n132, ZN => n1223);
   U104 : INV_X1 port map( A => n141, ZN => n1225);
   U105 : INV_X1 port map( A => n135, ZN => n1251);
   U106 : INV_X1 port map( A => n68, ZN => n1212);
   U107 : INV_X1 port map( A => n60, ZN => n1214);
   U108 : INV_X1 port map( A => n104, ZN => n1216);
   U109 : INV_X1 port map( A => n92, ZN => n1218);
   U110 : INV_X1 port map( A => n100, ZN => n1250);
   U111 : INV_X1 port map( A => SH(0), ZN => n1198);
   U112 : OAI221_X1 port map( B1 => n1232, B2 => n97, C1 => n1230, C2 => n98, A
                           => n159, ZN => n81);
   U113 : AOI22_X1 port map( A1 => A(20), A2 => n94, B1 => A(21), B2 => n95, ZN
                           => n159);
   U114 : OAI221_X1 port map( B1 => n1255, B2 => n1236, C1 => n1252, C2 => 
                           n1238, A => n158, ZN => n120);
   U115 : AOI22_X1 port map( A1 => A(23), A2 => n1254, B1 => A(22), B2 => n1253
                           , ZN => n158);
   U116 : OAI221_X1 port map( B1 => n1255, B2 => n1247, C1 => n1252, C2 => 
                           n1249, A => n171, ZN => n115);
   U117 : AOI22_X1 port map( A1 => A(29), A2 => n1254, B1 => A(28), B2 => n1253
                           , ZN => n171);
   U118 : OAI221_X1 port map( B1 => n97, B2 => n1234, C1 => n1233, C2 => n98, A
                           => n173, ZN => n72);
   U119 : INV_X1 port map( A => A(21), ZN => n1234);
   U120 : AOI22_X1 port map( A1 => A(22), A2 => n94, B1 => A(23), B2 => n95, ZN
                           => n173);
   U121 : OAI221_X1 port map( B1 => n1233, B2 => n97, C1 => n1232, C2 => n98, A
                           => n153, ZN => n77);
   U122 : AOI22_X1 port map( A1 => A(21), A2 => n94, B1 => A(22), B2 => n95, ZN
                           => n153);
   U123 : OAI221_X1 port map( B1 => n1255, B2 => n1238, C1 => n1252, C2 => 
                           n1240, A => n152, ZN => n118);
   U124 : AOI22_X1 port map( A1 => A(24), A2 => n1254, B1 => A(23), B2 => n1253
                           , ZN => n152);
   U125 : OAI221_X1 port map( B1 => n1255, B2 => n1240, C1 => n1252, C2 => 
                           n1241, A => n170, ZN => n116);
   U126 : AOI22_X1 port map( A1 => A(25), A2 => n1254, B1 => A(24), B2 => n1253
                           , ZN => n170);
   U127 : OAI221_X1 port map( B1 => n1255, B2 => n1241, C1 => n1252, C2 => 
                           n1243, A => n145, ZN => n113);
   U128 : AOI22_X1 port map( A1 => A(26), A2 => n1254, B1 => A(25), B2 => n1253
                           , ZN => n145);
   U129 : OAI221_X1 port map( B1 => n1255, B2 => n1235, C1 => n1252, C2 => 
                           n1236, A => n146, ZN => n67);
   U130 : INV_X1 port map( A => A(23), ZN => n1235);
   U131 : AOI22_X1 port map( A1 => A(22), A2 => n1254, B1 => A(21), B2 => n1253
                           , ZN => n146);
   U132 : OAI221_X1 port map( B1 => n1255, B2 => n1228, C1 => n1252, C2 => 
                           n1230, A => n154, ZN => n76);
   U133 : INV_X1 port map( A => A(17), ZN => n1228);
   U134 : AOI22_X1 port map( A1 => A(16), A2 => n1254, B1 => A(15), B2 => n1253
                           , ZN => n154);
   U135 : OAI221_X1 port map( B1 => n1255, B2 => n1230, C1 => n1232, C2 => 
                           n1252, A => n172, ZN => n71);
   U136 : AOI22_X1 port map( A1 => A(17), A2 => n1254, B1 => A(16), B2 => n1253
                           , ZN => n172);
   U137 : OAI221_X1 port map( B1 => n1255, B2 => n1232, C1 => n1252, C2 => 
                           n1233, A => n147, ZN => n65);
   U138 : AOI22_X1 port map( A1 => A(18), A2 => n1254, B1 => A(17), B2 => n1253
                           , ZN => n147);
   U139 : OAI221_X1 port map( B1 => n1255, B2 => n1246, C1 => n1252, C2 => 
                           n1247, A => n155, ZN => n117);
   U140 : AOI22_X1 port map( A1 => A(28), A2 => n1254, B1 => A(27), B2 => n1253
                           , ZN => n155);
   U141 : OAI221_X1 port map( B1 => n1255, B2 => n1243, C1 => n1252, C2 => 
                           n1246, A => n161, ZN => n119);
   U142 : AOI22_X1 port map( A1 => A(27), A2 => n1254, B1 => A(26), B2 => n1253
                           , ZN => n161);
   U143 : AOI221_X1 port map( B1 => n94, B2 => A(6), C1 => n95, C2 => A(7), A 
                           => n174, ZN => n85);
   U144 : OAI22_X1 port map( A1 => n1209, A2 => n97, B1 => n1208, B2 => n98, ZN
                           => n174);
   U145 : AOI221_X1 port map( B1 => n94, B2 => A(7), C1 => n95, C2 => A(8), A 
                           => n133, ZN => n82);
   U146 : OAI22_X1 port map( A1 => n1210, A2 => n97, B1 => n1209, B2 => n98, ZN
                           => n133);
   U147 : AOI221_X1 port map( B1 => n94, B2 => A(8), C1 => n95, C2 => A(9), A 
                           => n106, ZN => n78);
   U148 : OAI22_X1 port map( A1 => n1211, A2 => n97, B1 => n1210, B2 => n98, ZN
                           => n106);
   U149 : AOI221_X1 port map( B1 => n94, B2 => A(9), C1 => n95, C2 => A(10), A 
                           => n96, ZN => n73);
   U150 : OAI22_X1 port map( A1 => n1213, A2 => n97, B1 => n1211, B2 => n98, ZN
                           => n96);
   U151 : AOI221_X1 port map( B1 => n94, B2 => A(10), C1 => n95, C2 => A(11), A
                           => n165, ZN => n68);
   U152 : OAI22_X1 port map( A1 => n1215, A2 => n97, B1 => n1213, B2 => n98, ZN
                           => n165);
   U153 : AOI221_X1 port map( B1 => n94, B2 => A(11), C1 => n95, C2 => A(12), A
                           => n130, ZN => n60);
   U154 : OAI22_X1 port map( A1 => n1217, A2 => n97, B1 => n1215, B2 => n98, ZN
                           => n130);
   U155 : AOI221_X1 port map( B1 => n94, B2 => A(12), C1 => n95, C2 => A(13), A
                           => n162, ZN => n104);
   U156 : OAI22_X1 port map( A1 => n1219, A2 => n97, B1 => n1217, B2 => n98, ZN
                           => n162);
   U157 : AOI221_X1 port map( B1 => n94, B2 => A(13), C1 => n95, C2 => A(14), A
                           => n156, ZN => n92);
   U158 : OAI22_X1 port map( A1 => n1220, A2 => n97, B1 => n1219, B2 => n98, ZN
                           => n156);
   U159 : INV_X1 port map( A => A(12), ZN => n1220);
   U160 : AOI221_X1 port map( B1 => n94, B2 => A(14), C1 => n95, C2 => A(15), A
                           => n1222, ZN => n149);
   U161 : INV_X1 port map( A => n168, ZN => n1222);
   U162 : AOI22_X1 port map( A1 => A(13), A2 => n1254, B1 => A(12), B2 => n1253
                           , ZN => n168);
   U163 : AOI221_X1 port map( B1 => n94, B2 => A(15), C1 => n95, C2 => A(16), A
                           => n1224, ZN => n132);
   U164 : INV_X1 port map( A => n148, ZN => n1224);
   U165 : AOI22_X1 port map( A1 => A(14), A2 => n1254, B1 => A(13), B2 => n1253
                           , ZN => n148);
   U166 : AOI221_X1 port map( B1 => n94, B2 => A(16), C1 => n95, C2 => A(17), A
                           => n1226, ZN => n141);
   U167 : INV_X1 port map( A => n160, ZN => n1226);
   U168 : AOI22_X1 port map( A1 => A(15), A2 => n1254, B1 => A(14), B2 => n1253
                           , ZN => n160);
   U169 : OAI221_X1 port map( B1 => n82, B2 => n88, C1 => n127, C2 => n1203, A 
                           => n128, ZN => B_1_port);
   U170 : AOI222_X1 port map( A1 => n66, A2 => n1223, B1 => n1257, B2 => n129, 
                           C1 => n64, C2 => n1214, ZN => n128);
   U171 : OAI221_X1 port map( B1 => n1255, B2 => n1207, C1 => n1252, C2 => 
                           n1208, A => n131, ZN => n129);
   U172 : AOI22_X1 port map( A1 => A(2), A2 => n1254, B1 => A(1), B2 => n1253, 
                           ZN => n131);
   U173 : OAI221_X1 port map( B1 => n78, B2 => n88, C1 => n101, C2 => n1203, A 
                           => n102, ZN => B_2_port);
   U174 : AOI222_X1 port map( A1 => n66, A2 => n1225, B1 => n1257, B2 => n103, 
                           C1 => n64, C2 => n1216, ZN => n102);
   U175 : OAI221_X1 port map( B1 => n1255, B2 => n1208, C1 => n1252, C2 => 
                           n1209, A => n105, ZN => n103);
   U176 : AOI22_X1 port map( A1 => A(3), A2 => n1254, B1 => A(2), B2 => n1253, 
                           ZN => n105);
   U178 : OAI221_X1 port map( B1 => n73, B2 => n88, C1 => n89, C2 => n1203, A 
                           => n90, ZN => B_3_port);
   U179 : AOI222_X1 port map( A1 => n66, A2 => n76, B1 => n1257, B2 => n91, C1 
                           => n64, C2 => n1218, ZN => n90);
   U180 : OAI221_X1 port map( B1 => n1255, B2 => n1209, C1 => n1252, C2 => 
                           n1210, A => n93, ZN => n91);
   U181 : AOI22_X1 port map( A1 => A(4), A2 => n1254, B1 => A(3), B2 => n1253, 
                           ZN => n93);
   U182 : OAI221_X1 port map( B1 => n85, B2 => n88, C1 => n139, C2 => n1203, A 
                           => n163, ZN => B_0_port);
   U183 : AOI222_X1 port map( A1 => n66, A2 => n1221, B1 => n1257, B2 => n164, 
                           C1 => n64, C2 => n1212, ZN => n163);
   U184 : OAI221_X1 port map( B1 => n1255, B2 => n1206, C1 => n1252, C2 => 
                           n1207, A => n167, ZN => n164);
   U185 : INV_X1 port map( A => A(2), ZN => n1206);
   U186 : AOI22_X1 port map( A1 => A(1), A2 => n1254, B1 => A(0), B2 => n1253, 
                           ZN => n167);
   U187 : INV_X1 port map( A => A(5), ZN => n1209);
   U188 : INV_X1 port map( A => A(19), ZN => n1232);
   U189 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n135);
   U190 : INV_X1 port map( A => A(20), ZN => n1233);
   U191 : INV_X1 port map( A => A(31), ZN => n1249);
   U192 : INV_X1 port map( A => A(6), ZN => n1210);
   U193 : INV_X1 port map( A => A(4), ZN => n1208);
   U194 : INV_X1 port map( A => A(30), ZN => n1247);
   U195 : INV_X1 port map( A => A(18), ZN => n1230);
   U196 : INV_X1 port map( A => A(29), ZN => n1246);
   U197 : INV_X1 port map( A => A(26), ZN => n1240);
   U198 : INV_X1 port map( A => A(28), ZN => n1243);
   U199 : INV_X1 port map( A => A(27), ZN => n1241);
   U200 : INV_X1 port map( A => A(25), ZN => n1238);
   U201 : INV_X1 port map( A => A(24), ZN => n1236);
   U202 : INV_X1 port map( A => A(3), ZN => n1207);
   U203 : INV_X1 port map( A => A(8), ZN => n1213);
   U204 : INV_X1 port map( A => A(9), ZN => n1215);
   U205 : INV_X1 port map( A => A(10), ZN => n1217);
   U206 : INV_X1 port map( A => A(11), ZN => n1219);
   U207 : INV_X1 port map( A => A(7), ZN => n1211);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity adder_NBIT32_DW01_add_0_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end adder_NBIT32_DW01_add_0_DW01_add_1;

architecture SYN_rpl of adder_NBIT32_DW01_add_0_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1029 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1029, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity add4_NBIT32_DW01_add_0_DW01_add_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end add4_NBIT32_DW01_add_0_DW01_add_2;

architecture SYN_rpl of add4_NBIT32_DW01_add_0_DW01_add_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, SUM_31_port, n25, n26, n27, n28, 
      SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, 
      SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, 
      SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, 
      SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, SUM_11_port, 
      SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port, SUM_5_port, 
      SUM_4_port, SUM_3_port, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U30 : XOR2_X1 port map( A => A(30), B => n23, Z => SUM_30_port);
   U31 : XOR2_X1 port map( A => A(29), B => n22, Z => SUM_29_port);
   U32 : XOR2_X1 port map( A => A(28), B => n21, Z => SUM_28_port);
   U33 : XOR2_X1 port map( A => A(27), B => n20, Z => SUM_27_port);
   U34 : XOR2_X1 port map( A => A(26), B => n19, Z => SUM_26_port);
   U35 : XOR2_X1 port map( A => A(25), B => n18, Z => SUM_25_port);
   U36 : XOR2_X1 port map( A => A(24), B => n17, Z => SUM_24_port);
   U37 : XOR2_X1 port map( A => A(23), B => n16, Z => SUM_23_port);
   U38 : XOR2_X1 port map( A => A(22), B => n15, Z => SUM_22_port);
   U39 : XOR2_X1 port map( A => A(21), B => n14, Z => SUM_21_port);
   U40 : XOR2_X1 port map( A => A(20), B => n13, Z => SUM_20_port);
   U41 : XOR2_X1 port map( A => A(19), B => n12, Z => SUM_19_port);
   U42 : XOR2_X1 port map( A => A(18), B => n11, Z => SUM_18_port);
   U43 : XOR2_X1 port map( A => A(17), B => n10, Z => SUM_17_port);
   U44 : XOR2_X1 port map( A => A(16), B => n9, Z => SUM_16_port);
   U45 : XOR2_X1 port map( A => A(15), B => n8, Z => SUM_15_port);
   U46 : XOR2_X1 port map( A => A(14), B => n7, Z => SUM_14_port);
   U47 : XOR2_X1 port map( A => A(13), B => n6, Z => SUM_13_port);
   U48 : XOR2_X1 port map( A => A(12), B => n28, Z => SUM_12_port);
   U49 : XOR2_X1 port map( A => A(11), B => n5, Z => SUM_11_port);
   U50 : XOR2_X1 port map( A => A(10), B => n27, Z => SUM_10_port);
   U51 : XOR2_X1 port map( A => A(9), B => n4, Z => SUM_9_port);
   U52 : XOR2_X1 port map( A => A(8), B => n26, Z => SUM_8_port);
   U53 : XOR2_X1 port map( A => A(7), B => n3, Z => SUM_7_port);
   U54 : XOR2_X1 port map( A => A(6), B => n2, Z => SUM_6_port);
   U55 : XOR2_X1 port map( A => A(5), B => n1, Z => SUM_5_port);
   U56 : XOR2_X1 port map( A => A(4), B => n25, Z => SUM_4_port);
   U57 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U1 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U2 : NAND2_X1 port map( A1 => A(30), A2 => n23, ZN => n57);
   U3 : AND2_X1 port map( A1 => A(29), A2 => n22, ZN => n23);
   U4 : AND2_X1 port map( A1 => A(4), A2 => n25, ZN => n1);
   U5 : AND2_X1 port map( A1 => A(5), A2 => n1, ZN => n2);
   U6 : AND2_X1 port map( A1 => A(6), A2 => n2, ZN => n3);
   U7 : AND2_X1 port map( A1 => A(7), A2 => n3, ZN => n26);
   U8 : AND2_X1 port map( A1 => A(8), A2 => n26, ZN => n4);
   U9 : AND2_X1 port map( A1 => A(9), A2 => n4, ZN => n27);
   U10 : AND2_X1 port map( A1 => A(10), A2 => n27, ZN => n5);
   U11 : AND2_X1 port map( A1 => A(11), A2 => n5, ZN => n28);
   U12 : AND2_X1 port map( A1 => A(12), A2 => n28, ZN => n6);
   U13 : AND2_X1 port map( A1 => A(13), A2 => n6, ZN => n7);
   U14 : AND2_X1 port map( A1 => A(14), A2 => n7, ZN => n8);
   U15 : AND2_X1 port map( A1 => A(15), A2 => n8, ZN => n9);
   U16 : AND2_X1 port map( A1 => A(16), A2 => n9, ZN => n10);
   U17 : AND2_X1 port map( A1 => A(17), A2 => n10, ZN => n11);
   U18 : AND2_X1 port map( A1 => A(18), A2 => n11, ZN => n12);
   U19 : AND2_X1 port map( A1 => A(19), A2 => n12, ZN => n13);
   U20 : AND2_X1 port map( A1 => A(20), A2 => n13, ZN => n14);
   U21 : AND2_X1 port map( A1 => A(21), A2 => n14, ZN => n15);
   U22 : AND2_X1 port map( A1 => A(22), A2 => n15, ZN => n16);
   U23 : AND2_X1 port map( A1 => A(23), A2 => n16, ZN => n17);
   U24 : AND2_X1 port map( A1 => A(24), A2 => n17, ZN => n18);
   U25 : AND2_X1 port map( A1 => A(25), A2 => n18, ZN => n19);
   U26 : AND2_X1 port map( A1 => A(26), A2 => n19, ZN => n20);
   U27 : AND2_X1 port map( A1 => A(27), A2 => n20, ZN => n21);
   U28 : AND2_X1 port map( A1 => A(28), A2 => n21, ZN => n22);
   U29 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n25);
   U58 : INV_X1 port map( A => A(2), ZN => SUM_2_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity is_zero_NBIT32 is

   port( A : in std_logic_vector (31 downto 0);  BEQZ_OR_BNEZ, EN : in 
         std_logic;  res : out std_logic);

end is_zero_NBIT32;

architecture SYN_beh of is_zero_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U3 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n8);
   U4 : NOR4_X1 port map( A1 => n13, A2 => A(8), A3 => BEQZ_OR_BNEZ, A4 => A(9)
                           , ZN => n12);
   U5 : OR2_X1 port map( A1 => A(7), A2 => A(6), ZN => n13);
   U6 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), ZN
                           => n7);
   U7 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n11);
   U8 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n6);
   U9 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), ZN
                           => n10);
   U10 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), 
                           ZN => n5);
   U11 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n9);
   U12 : OAI21_X1 port map( B1 => n3, B2 => n4, A => EN, ZN => n2);
   U13 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n3
                           );
   U14 : NAND4_X1 port map( A1 => n5, A2 => n6, A3 => n7, A4 => n8, ZN => n4);
   U15 : INV_X1 port map( A => n2, ZN => res);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32 is

   port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end ALU_N32;

architecture SYN_BEHAVIOR of ALU_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ALU_N32_DW02_mult_0
      port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_N32_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component ALU_N32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component ALU_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component ALU_N32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal tmp_sub_31_port, tmp_sub_30_port, tmp_sub_29_port, tmp_sub_28_port, 
      tmp_sub_27_port, tmp_sub_26_port, tmp_sub_25_port, tmp_sub_24_port, 
      tmp_sub_23_port, tmp_sub_22_port, tmp_sub_21_port, tmp_sub_20_port, 
      tmp_sub_19_port, tmp_sub_18_port, tmp_sub_17_port, tmp_sub_16_port, 
      tmp_sub_15_port, tmp_sub_14_port, tmp_sub_13_port, tmp_sub_12_port, 
      tmp_sub_11_port, tmp_sub_10_port, tmp_sub_9_port, tmp_sub_8_port, 
      tmp_sub_7_port, tmp_sub_6_port, tmp_sub_5_port, tmp_sub_4_port, 
      tmp_sub_3_port, tmp_sub_2_port, tmp_sub_1_port, tmp_sub_0_port, N78, N79,
      N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94
      , N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107
      , N108, N109, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
      N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, 
      N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, 
      N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, 
      N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, 
      N332, N333, n6, n7, n8, n9, n10, n81_port, n82_port, n83_port, n84_port, 
      n85_port, n86_port, n87_port, n88_port, n89_port, n90_port, n91_port, 
      n92_port, n93_port, n94_port, n95_port, n96_port, n97_port, n98_port, 
      n99_port, n100_port, n101_port, n102_port, n103_port, n104_port, 
      n105_port, n106_port, n107_port, n108_port, n109_port, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142_port, n143_port, n144_port, n145_port,
      n146_port, n147_port, n148_port, n149_port, n150_port, n151_port, 
      n152_port, n153_port, n154_port, n155_port, n156_port, n157_port, 
      n158_port, n159_port, n160_port, n161_port, n162_port, n163_port, 
      n164_port, n165_port, n166_port, n167_port, n168_port, n169_port, 
      n170_port, n171_port, n172_port, n173_port, n174, n175, n176, n177, n178,
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
      n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, 
      n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, 
      n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, 
      n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, 
      n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
      n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, 
      n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, 
      n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, 
      n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, 
      n2468, n2469, n2470, n2471, n2472, n2473, n_1064, n_1065 : std_logic;

begin
   
   n6 <= '0';
   n7 <= '0';
   n8 <= '1';
   n9 <= '0';
   n10 <= '0';
   U293 : NAND3_X1 port map( A1 => n243, A2 => n244, A3 => n245, ZN => 
                           OUTALU(0));
   U294 : OAI33_X1 port map( A1 => n2410, A2 => DATA2(0), A3 => n247, B1 => 
                           n248, B2 => n249, B3 => n2470, ZN => n246);
   U295 : NAND3_X1 port map( A1 => n2472, A2 => n2470, A3 => FUNC(1), ZN => 
                           n247);
   sra_42 : ALU_N32_DW_sra_0 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), SH(4) => DATA2(4), 
                           SH(3) => DATA2(3), SH(2) => DATA2(2), SH(1) => 
                           DATA2(1), SH(0) => DATA2(0), SH_TC => n9, B(31) => 
                           N333, B(30) => N332, B(29) => N331, B(28) => N330, 
                           B(27) => N329, B(26) => N328, B(25) => N327, B(24) 
                           => N326, B(23) => N325, B(22) => N324, B(21) => N323
                           , B(20) => N322, B(19) => N321, B(18) => N320, B(17)
                           => N319, B(16) => N318, B(15) => N317, B(14) => N316
                           , B(13) => N315, B(12) => N314, B(11) => N313, B(10)
                           => N312, B(9) => N311, B(8) => N310, B(7) => N309, 
                           B(6) => N308, B(5) => N307, B(4) => N306, B(3) => 
                           N305, B(2) => N304, B(1) => N303, B(0) => N302);
   sll_41 : ALU_N32_DW01_ash_0 port map( A(31) => DATA1(31), A(30) => DATA1(30)
                           , A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), DATA_TC => n10, SH(4)
                           => DATA2(4), SH(3) => DATA2(3), SH(2) => DATA2(2), 
                           SH(1) => DATA2(1), SH(0) => DATA2(0), SH_TC => n10, 
                           B(31) => N301, B(30) => N300, B(29) => N299, B(28) 
                           => N298, B(27) => N297, B(26) => N296, B(25) => N295
                           , B(24) => N294, B(23) => N293, B(22) => N292, B(21)
                           => N291, B(20) => N290, B(19) => N289, B(18) => N288
                           , B(17) => N287, B(16) => N286, B(15) => N285, B(14)
                           => N284, B(13) => N283, B(12) => N282, B(11) => N281
                           , B(10) => N280, B(9) => N279, B(8) => N278, B(7) =>
                           N277, B(6) => N276, B(5) => N275, B(4) => N274, B(3)
                           => N273, B(2) => N272, B(1) => N271, B(0) => N270);
   add_35 : ALU_N32_DW01_add_0 port map( A(31) => DATA1(31), A(30) => DATA1(30)
                           , A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , CI => n6, SUM(31) => N109, SUM(30) => N108, 
                           SUM(29) => N107, SUM(28) => N106, SUM(27) => N105, 
                           SUM(26) => N104, SUM(25) => N103, SUM(24) => N102, 
                           SUM(23) => N101, SUM(22) => N100, SUM(21) => N99, 
                           SUM(20) => N98, SUM(19) => N97, SUM(18) => N96, 
                           SUM(17) => N95, SUM(16) => N94, SUM(15) => N93, 
                           SUM(14) => N92, SUM(13) => N91, SUM(12) => N90, 
                           SUM(11) => N89, SUM(10) => N88, SUM(9) => N87, 
                           SUM(8) => N86, SUM(7) => N85, SUM(6) => N84, SUM(5) 
                           => N83, SUM(4) => N82, SUM(3) => N81, SUM(2) => N80,
                           SUM(1) => N79, SUM(0) => N78, CO => n_1064);
   r62 : ALU_N32_DW01_sub_0 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , CI => n7, DIFF(31) => tmp_sub_31_port, DIFF(30) =>
                           tmp_sub_30_port, DIFF(29) => tmp_sub_29_port, 
                           DIFF(28) => tmp_sub_28_port, DIFF(27) => 
                           tmp_sub_27_port, DIFF(26) => tmp_sub_26_port, 
                           DIFF(25) => tmp_sub_25_port, DIFF(24) => 
                           tmp_sub_24_port, DIFF(23) => tmp_sub_23_port, 
                           DIFF(22) => tmp_sub_22_port, DIFF(21) => 
                           tmp_sub_21_port, DIFF(20) => tmp_sub_20_port, 
                           DIFF(19) => tmp_sub_19_port, DIFF(18) => 
                           tmp_sub_18_port, DIFF(17) => tmp_sub_17_port, 
                           DIFF(16) => tmp_sub_16_port, DIFF(15) => 
                           tmp_sub_15_port, DIFF(14) => tmp_sub_14_port, 
                           DIFF(13) => tmp_sub_13_port, DIFF(12) => 
                           tmp_sub_12_port, DIFF(11) => tmp_sub_11_port, 
                           DIFF(10) => tmp_sub_10_port, DIFF(9) => 
                           tmp_sub_9_port, DIFF(8) => tmp_sub_8_port, DIFF(7) 
                           => tmp_sub_7_port, DIFF(6) => tmp_sub_6_port, 
                           DIFF(5) => tmp_sub_5_port, DIFF(4) => tmp_sub_4_port
                           , DIFF(3) => tmp_sub_3_port, DIFF(2) => 
                           tmp_sub_2_port, DIFF(1) => tmp_sub_1_port, DIFF(0) 
                           => tmp_sub_0_port, CO => n_1065);
   mult_37 : ALU_N32_DW02_mult_0 port map( A(15) => DATA1(15), A(14) => 
                           DATA1(14), A(13) => DATA1(13), A(12) => DATA1(12), 
                           A(11) => DATA1(11), A(10) => DATA1(10), A(9) => 
                           DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7), A(6) 
                           => DATA1(6), A(5) => DATA1(5), A(4) => DATA1(4), 
                           A(3) => DATA1(3), A(2) => DATA1(2), A(1) => DATA1(1)
                           , A(0) => DATA1(0), B(15) => DATA2(15), B(14) => 
                           DATA2(14), B(13) => DATA2(13), B(12) => DATA2(12), 
                           B(11) => DATA2(11), B(10) => DATA2(10), B(9) => 
                           DATA2(9), B(8) => DATA2(8), B(7) => DATA2(7), B(6) 
                           => DATA2(6), B(5) => DATA2(5), B(4) => DATA2(4), 
                           B(3) => DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1)
                           , B(0) => DATA2(0), TC => n8, PRODUCT(31) => N173, 
                           PRODUCT(30) => N172, PRODUCT(29) => N171, 
                           PRODUCT(28) => N170, PRODUCT(27) => N169, 
                           PRODUCT(26) => N168, PRODUCT(25) => N167, 
                           PRODUCT(24) => N166, PRODUCT(23) => N165, 
                           PRODUCT(22) => N164, PRODUCT(21) => N163, 
                           PRODUCT(20) => N162, PRODUCT(19) => N161, 
                           PRODUCT(18) => N160, PRODUCT(17) => N159, 
                           PRODUCT(16) => N158, PRODUCT(15) => N157, 
                           PRODUCT(14) => N156, PRODUCT(13) => N155, 
                           PRODUCT(12) => N154, PRODUCT(11) => N153, 
                           PRODUCT(10) => N152, PRODUCT(9) => N151, PRODUCT(8) 
                           => N150, PRODUCT(7) => N149, PRODUCT(6) => N148, 
                           PRODUCT(5) => N147, PRODUCT(4) => N146, PRODUCT(3) 
                           => N145, PRODUCT(2) => N144, PRODUCT(1) => N143, 
                           PRODUCT(0) => N142);
   U4 : BUF_X1 port map( A => n2469, Z => n2375);
   U5 : BUF_X1 port map( A => n2469, Z => n2374);
   U6 : BUF_X1 port map( A => n90_port, Z => n2384);
   U7 : BUF_X1 port map( A => n84_port, Z => n2399);
   U10 : BUF_X1 port map( A => n83_port, Z => n2403);
   U12 : BUF_X1 port map( A => n89_port, Z => n2391);
   U13 : BUF_X1 port map( A => n88_port, Z => n2392);
   U14 : BUF_X1 port map( A => n91_port, Z => n2380);
   U15 : BUF_X1 port map( A => n92_port, Z => n2376);
   U16 : BUF_X1 port map( A => n2374, Z => n2372);
   U17 : BUF_X1 port map( A => n2374, Z => n2371);
   U18 : BUF_X1 port map( A => n2375, Z => n2368);
   U19 : BUF_X1 port map( A => n2375, Z => n2369);
   U20 : BUF_X1 port map( A => n2375, Z => n2370);
   U21 : BUF_X1 port map( A => n2374, Z => n2373);
   U22 : BUF_X1 port map( A => n2384, Z => n2385);
   U23 : BUF_X1 port map( A => n2384, Z => n2386);
   U24 : BUF_X1 port map( A => n2384, Z => n2387);
   U25 : NOR4_X1 port map( A1 => tmp_sub_9_port, A2 => tmp_sub_8_port, A3 => 
                           tmp_sub_7_port, A4 => tmp_sub_6_port, ZN => n260);
   U26 : NOR4_X1 port map( A1 => tmp_sub_22_port, A2 => tmp_sub_21_port, A3 => 
                           tmp_sub_20_port, A4 => tmp_sub_1_port, ZN => n256);
   U27 : NOR4_X1 port map( A1 => tmp_sub_5_port, A2 => tmp_sub_4_port, A3 => 
                           tmp_sub_3_port, A4 => tmp_sub_30_port, ZN => n259);
   U28 : NOR4_X1 port map( A1 => tmp_sub_19_port, A2 => tmp_sub_18_port, A3 => 
                           tmp_sub_17_port, A4 => tmp_sub_16_port, ZN => n255);
   U29 : NOR4_X1 port map( A1 => tmp_sub_2_port, A2 => tmp_sub_29_port, A3 => 
                           tmp_sub_28_port, A4 => tmp_sub_27_port, ZN => n258);
   U30 : NOR4_X1 port map( A1 => tmp_sub_15_port, A2 => tmp_sub_14_port, A3 => 
                           tmp_sub_13_port, A4 => tmp_sub_12_port, ZN => n254);
   U31 : NOR4_X1 port map( A1 => tmp_sub_26_port, A2 => tmp_sub_25_port, A3 => 
                           tmp_sub_24_port, A4 => tmp_sub_23_port, ZN => n257);
   U32 : NAND2_X1 port map( A1 => n188, A2 => n189, ZN => OUTALU(1));
   U33 : AOI221_X1 port map( B1 => N303, B2 => n2400, C1 => N271, C2 => n2397, 
                           A => n190, ZN => n189);
   U34 : AOI222_X1 port map( A1 => N79, A2 => n2385, B1 => N143, B2 => n2381, 
                           C1 => tmp_sub_1_port, C2 => n2377, ZN => n188);
   U35 : NAND2_X1 port map( A1 => n133, A2 => n134, ZN => OUTALU(2));
   U36 : AOI221_X1 port map( B1 => N304, B2 => n2401, C1 => N272, C2 => n2396, 
                           A => n135, ZN => n134);
   U37 : AOI222_X1 port map( A1 => N80, A2 => n2386, B1 => N144, B2 => n2382, 
                           C1 => tmp_sub_2_port, C2 => n2378, ZN => n133);
   U38 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => OUTALU(3));
   U39 : AOI221_X1 port map( B1 => N305, B2 => n2402, C1 => N273, C2 => n2396, 
                           A => n120, ZN => n119);
   U40 : AOI222_X1 port map( A1 => N81, A2 => n2387, B1 => N145, B2 => n2383, 
                           C1 => tmp_sub_3_port, C2 => n2379, ZN => n118);
   U41 : NAND2_X1 port map( A1 => n113, A2 => n114, ZN => OUTALU(4));
   U42 : AOI221_X1 port map( B1 => N306, B2 => n2402, C1 => N274, C2 => n2396, 
                           A => n115, ZN => n114);
   U43 : AOI222_X1 port map( A1 => N82, A2 => n2387, B1 => N146, B2 => n2383, 
                           C1 => tmp_sub_4_port, C2 => n2379, ZN => n113);
   U44 : NAND2_X1 port map( A1 => n108_port, A2 => n109_port, ZN => OUTALU(5));
   U45 : AOI221_X1 port map( B1 => N307, B2 => n2402, C1 => N275, C2 => n2396, 
                           A => n110, ZN => n109_port);
   U46 : AOI222_X1 port map( A1 => N83, A2 => n2387, B1 => N147, B2 => n2383, 
                           C1 => tmp_sub_5_port, C2 => n2379, ZN => n108_port);
   U47 : NAND2_X1 port map( A1 => n103_port, A2 => n104_port, ZN => OUTALU(6));
   U48 : AOI221_X1 port map( B1 => N308, B2 => n2402, C1 => N276, C2 => n2396, 
                           A => n105_port, ZN => n104_port);
   U49 : AOI222_X1 port map( A1 => N84, A2 => n2387, B1 => N148, B2 => n2383, 
                           C1 => tmp_sub_6_port, C2 => n2379, ZN => n103_port);
   U50 : NAND2_X1 port map( A1 => n98_port, A2 => n99_port, ZN => OUTALU(7));
   U51 : AOI221_X1 port map( B1 => N309, B2 => n2402, C1 => N277, C2 => n2396, 
                           A => n100_port, ZN => n99_port);
   U52 : AOI222_X1 port map( A1 => N85, A2 => n2387, B1 => N149, B2 => n2383, 
                           C1 => tmp_sub_7_port, C2 => n2379, ZN => n98_port);
   U53 : NAND2_X1 port map( A1 => n93_port, A2 => n94_port, ZN => OUTALU(8));
   U54 : AOI221_X1 port map( B1 => N310, B2 => n2402, C1 => N278, C2 => n2396, 
                           A => n95_port, ZN => n94_port);
   U55 : AOI222_X1 port map( A1 => N86, A2 => n2387, B1 => N150, B2 => n2383, 
                           C1 => tmp_sub_8_port, C2 => n2379, ZN => n93_port);
   U56 : NAND2_X1 port map( A1 => n81_port, A2 => n82_port, ZN => OUTALU(9));
   U57 : AOI221_X1 port map( B1 => N311, B2 => n2402, C1 => N279, C2 => n2396, 
                           A => n85_port, ZN => n82_port);
   U58 : AOI222_X1 port map( A1 => N87, A2 => n2387, B1 => N151, B2 => n2383, 
                           C1 => tmp_sub_9_port, C2 => n2379, ZN => n81_port);
   U59 : NAND2_X1 port map( A1 => n238, A2 => n239, ZN => OUTALU(10));
   U60 : AOI221_X1 port map( B1 => N312, B2 => n2400, C1 => N280, C2 => n2398, 
                           A => n240, ZN => n239);
   U61 : AOI222_X1 port map( A1 => N88, A2 => n2385, B1 => N152, B2 => n2381, 
                           C1 => tmp_sub_10_port, C2 => n2377, ZN => n238);
   U62 : NAND2_X1 port map( A1 => n233, A2 => n234, ZN => OUTALU(11));
   U63 : AOI221_X1 port map( B1 => N313, B2 => n2400, C1 => N281, C2 => n2398, 
                           A => n235, ZN => n234);
   U64 : AOI222_X1 port map( A1 => N89, A2 => n2385, B1 => N153, B2 => n2381, 
                           C1 => tmp_sub_11_port, C2 => n2377, ZN => n233);
   U65 : NAND2_X1 port map( A1 => n228, A2 => n229, ZN => OUTALU(12));
   U66 : AOI221_X1 port map( B1 => N314, B2 => n2400, C1 => N282, C2 => n2398, 
                           A => n230, ZN => n229);
   U67 : AOI222_X1 port map( A1 => N90, A2 => n2385, B1 => N154, B2 => n2381, 
                           C1 => tmp_sub_12_port, C2 => n2377, ZN => n228);
   U68 : NAND2_X1 port map( A1 => n223, A2 => n224, ZN => OUTALU(13));
   U69 : AOI221_X1 port map( B1 => N315, B2 => n2400, C1 => N283, C2 => n2398, 
                           A => n225, ZN => n224);
   U70 : AOI222_X1 port map( A1 => N91, A2 => n2385, B1 => N155, B2 => n2381, 
                           C1 => tmp_sub_13_port, C2 => n2377, ZN => n223);
   U71 : NAND2_X1 port map( A1 => n218, A2 => n219, ZN => OUTALU(14));
   U72 : AOI221_X1 port map( B1 => N316, B2 => n2400, C1 => N284, C2 => n2398, 
                           A => n220, ZN => n219);
   U73 : AOI222_X1 port map( A1 => N92, A2 => n2385, B1 => N156, B2 => n2381, 
                           C1 => tmp_sub_14_port, C2 => n2377, ZN => n218);
   U74 : NAND2_X1 port map( A1 => n213, A2 => n214, ZN => OUTALU(15));
   U75 : AOI221_X1 port map( B1 => N317, B2 => n2400, C1 => N285, C2 => n2398, 
                           A => n215, ZN => n214);
   U76 : AOI222_X1 port map( A1 => N93, A2 => n2385, B1 => N157, B2 => n2381, 
                           C1 => tmp_sub_15_port, C2 => n2377, ZN => n213);
   U77 : NAND2_X1 port map( A1 => n208, A2 => n209, ZN => OUTALU(16));
   U78 : AOI221_X1 port map( B1 => N318, B2 => n2400, C1 => N286, C2 => n2398, 
                           A => n210, ZN => n209);
   U79 : AOI222_X1 port map( A1 => N94, A2 => n2385, B1 => N158, B2 => n2381, 
                           C1 => tmp_sub_16_port, C2 => n2377, ZN => n208);
   U80 : NAND2_X1 port map( A1 => n203, A2 => n204, ZN => OUTALU(17));
   U81 : AOI221_X1 port map( B1 => N319, B2 => n2400, C1 => N287, C2 => n2397, 
                           A => n205, ZN => n204);
   U82 : AOI222_X1 port map( A1 => N95, A2 => n2385, B1 => N159, B2 => n2381, 
                           C1 => tmp_sub_17_port, C2 => n2377, ZN => n203);
   U83 : NAND2_X1 port map( A1 => n198, A2 => n199, ZN => OUTALU(18));
   U84 : AOI221_X1 port map( B1 => N320, B2 => n2400, C1 => N288, C2 => n2397, 
                           A => n200, ZN => n199);
   U85 : AOI222_X1 port map( A1 => N96, A2 => n2385, B1 => N160, B2 => n2381, 
                           C1 => tmp_sub_18_port, C2 => n2377, ZN => n198);
   U86 : NAND2_X1 port map( A1 => n193, A2 => n194, ZN => OUTALU(19));
   U87 : AOI221_X1 port map( B1 => N321, B2 => n2400, C1 => N289, C2 => n2397, 
                           A => n195, ZN => n194);
   U88 : AOI222_X1 port map( A1 => N97, A2 => n2385, B1 => N161, B2 => n2381, 
                           C1 => tmp_sub_19_port, C2 => n2377, ZN => n193);
   U89 : NAND2_X1 port map( A1 => n183, A2 => n184, ZN => OUTALU(20));
   U90 : AOI221_X1 port map( B1 => N322, B2 => n2401, C1 => N290, C2 => n2397, 
                           A => n185, ZN => n184);
   U91 : AOI222_X1 port map( A1 => N98, A2 => n2386, B1 => N162, B2 => n2382, 
                           C1 => tmp_sub_20_port, C2 => n2378, ZN => n183);
   U92 : NAND2_X1 port map( A1 => n178, A2 => n179, ZN => OUTALU(21));
   U93 : AOI221_X1 port map( B1 => N323, B2 => n2401, C1 => N291, C2 => n2397, 
                           A => n180, ZN => n179);
   U94 : AOI222_X1 port map( A1 => N99, A2 => n2386, B1 => N163, B2 => n2382, 
                           C1 => tmp_sub_21_port, C2 => n2378, ZN => n178);
   U95 : NAND2_X1 port map( A1 => n173_port, A2 => n174, ZN => OUTALU(22));
   U96 : AOI221_X1 port map( B1 => N324, B2 => n2401, C1 => N292, C2 => n2397, 
                           A => n175, ZN => n174);
   U97 : AOI222_X1 port map( A1 => N100, A2 => n2386, B1 => N164, B2 => n2382, 
                           C1 => tmp_sub_22_port, C2 => n2378, ZN => n173_port)
                           ;
   U98 : NAND2_X1 port map( A1 => n168_port, A2 => n169_port, ZN => OUTALU(23))
                           ;
   U99 : AOI221_X1 port map( B1 => N325, B2 => n2401, C1 => N293, C2 => n2397, 
                           A => n170_port, ZN => n169_port);
   U100 : AOI222_X1 port map( A1 => N101, A2 => n2386, B1 => N165, B2 => n2382,
                           C1 => tmp_sub_23_port, C2 => n2378, ZN => n168_port)
                           ;
   U101 : NAND2_X1 port map( A1 => n163_port, A2 => n164_port, ZN => OUTALU(24)
                           );
   U102 : AOI221_X1 port map( B1 => N326, B2 => n2401, C1 => N294, C2 => n2397,
                           A => n165_port, ZN => n164_port);
   U103 : AOI222_X1 port map( A1 => N102, A2 => n2386, B1 => N166, B2 => n2382,
                           C1 => tmp_sub_24_port, C2 => n2378, ZN => n163_port)
                           ;
   U104 : NAND2_X1 port map( A1 => n158_port, A2 => n159_port, ZN => OUTALU(25)
                           );
   U105 : AOI221_X1 port map( B1 => N327, B2 => n2401, C1 => N295, C2 => n2397,
                           A => n160_port, ZN => n159_port);
   U106 : AOI222_X1 port map( A1 => N103, A2 => n2386, B1 => N167, B2 => n2382,
                           C1 => tmp_sub_25_port, C2 => n2378, ZN => n158_port)
                           ;
   U107 : NAND2_X1 port map( A1 => n153_port, A2 => n154_port, ZN => OUTALU(26)
                           );
   U108 : AOI221_X1 port map( B1 => N328, B2 => n2401, C1 => N296, C2 => n2397,
                           A => n155_port, ZN => n154_port);
   U109 : AOI222_X1 port map( A1 => N104, A2 => n2386, B1 => N168, B2 => n2382,
                           C1 => tmp_sub_26_port, C2 => n2378, ZN => n153_port)
                           ;
   U110 : NAND2_X1 port map( A1 => n148_port, A2 => n149_port, ZN => OUTALU(27)
                           );
   U111 : AOI221_X1 port map( B1 => N329, B2 => n2401, C1 => N297, C2 => n2397,
                           A => n150_port, ZN => n149_port);
   U112 : AOI222_X1 port map( A1 => N105, A2 => n2386, B1 => N169, B2 => n2382,
                           C1 => tmp_sub_27_port, C2 => n2378, ZN => n148_port)
                           ;
   U113 : NAND2_X1 port map( A1 => n143_port, A2 => n144_port, ZN => OUTALU(28)
                           );
   U114 : AOI221_X1 port map( B1 => N330, B2 => n2401, C1 => N298, C2 => n2396,
                           A => n145_port, ZN => n144_port);
   U115 : AOI222_X1 port map( A1 => N106, A2 => n2386, B1 => N170, B2 => n2382,
                           C1 => tmp_sub_28_port, C2 => n2378, ZN => n143_port)
                           ;
   U116 : NAND2_X1 port map( A1 => n138, A2 => n139, ZN => OUTALU(29));
   U117 : AOI221_X1 port map( B1 => N331, B2 => n2401, C1 => N299, C2 => n2396,
                           A => n140, ZN => n139);
   U118 : AOI222_X1 port map( A1 => N107, A2 => n2386, B1 => N171, B2 => n2382,
                           C1 => tmp_sub_29_port, C2 => n2378, ZN => n138);
   U119 : NAND2_X1 port map( A1 => n128, A2 => n129, ZN => OUTALU(30));
   U120 : AOI221_X1 port map( B1 => N332, B2 => n2401, C1 => N300, C2 => n2396,
                           A => n130, ZN => n129);
   U121 : AOI222_X1 port map( A1 => N108, A2 => n2386, B1 => N172, B2 => n2382,
                           C1 => tmp_sub_30_port, C2 => n2378, ZN => n128);
   U122 : AOI22_X1 port map( A1 => tmp_sub_0_port, A2 => n2377, B1 => N78, B2 
                           => n2385, ZN => n243);
   U123 : AOI22_X1 port map( A1 => N270, A2 => n2398, B1 => N142, B2 => n2381, 
                           ZN => n244);
   U124 : AOI221_X1 port map( B1 => DATA2(0), B2 => n2409, C1 => N302, C2 => 
                           n2400, A => n246, ZN => n245);
   U125 : AND3_X1 port map( A1 => n2473, A2 => n2472, A3 => n262, ZN => 
                           n90_port);
   U126 : INV_X1 port map( A => n247, ZN => n2469);
   U127 : BUF_X1 port map( A => n2399, Z => n2397);
   U128 : BUF_X1 port map( A => n2399, Z => n2396);
   U129 : BUF_X1 port map( A => n2403, Z => n2401);
   U130 : BUF_X1 port map( A => n2391, Z => n2388);
   U131 : BUF_X1 port map( A => n2391, Z => n2389);
   U132 : BUF_X1 port map( A => n2380, Z => n2381);
   U133 : BUF_X1 port map( A => n2380, Z => n2382);
   U134 : BUF_X1 port map( A => n2376, Z => n2377);
   U135 : BUF_X1 port map( A => n2376, Z => n2378);
   U136 : BUF_X1 port map( A => n2403, Z => n2400);
   U137 : BUF_X1 port map( A => n2392, Z => n2393);
   U138 : BUF_X1 port map( A => n2392, Z => n2394);
   U139 : BUF_X1 port map( A => n2399, Z => n2398);
   U140 : BUF_X1 port map( A => n2391, Z => n2390);
   U141 : BUF_X1 port map( A => n2380, Z => n2383);
   U142 : BUF_X1 port map( A => n2376, Z => n2379);
   U143 : BUF_X1 port map( A => n2392, Z => n2395);
   U144 : BUF_X1 port map( A => n2403, Z => n2402);
   U145 : NAND2_X1 port map( A1 => n2472, A2 => n2471, ZN => n248);
   U146 : AOI22_X1 port map( A1 => n250, A2 => n2408, B1 => tmp_sub_31_port, B2
                           => FUNC(3), ZN => n249);
   U147 : INV_X1 port map( A => tmp_sub_31_port, ZN => n2408);
   U148 : OAI22_X1 port map( A1 => n191, A2 => n2411, B1 => n2404, B2 => n192, 
                           ZN => n190);
   U149 : NAND2_X1 port map( A1 => n2372, A2 => n2411, ZN => n192);
   U150 : INV_X1 port map( A => DATA1(1), ZN => n2411);
   U151 : AOI221_X1 port map( B1 => DATA2(1), B2 => n2394, C1 => n2369, C2 => 
                           n2404, A => n2388, ZN => n191);
   U152 : OAI22_X1 port map( A1 => n136, A2 => n2405, B1 => n2412, B2 => n137, 
                           ZN => n135);
   U153 : NAND2_X1 port map( A1 => n2371, A2 => n2405, ZN => n137);
   U154 : AOI221_X1 port map( B1 => DATA1(2), B2 => n2393, C1 => n2370, C2 => 
                           n2412, A => n2389, ZN => n136);
   U155 : INV_X1 port map( A => DATA1(2), ZN => n2412);
   U156 : OAI22_X1 port map( A1 => n121, A2 => n2413, B1 => n2406, B2 => n122, 
                           ZN => n120);
   U157 : NAND2_X1 port map( A1 => n2371, A2 => n2413, ZN => n122);
   U158 : INV_X1 port map( A => DATA1(3), ZN => n2413);
   U159 : AOI221_X1 port map( B1 => DATA2(3), B2 => n2393, C1 => n2370, C2 => 
                           n2406, A => n2390, ZN => n121);
   U160 : OAI22_X1 port map( A1 => n116, A2 => n2407, B1 => n2414, B2 => n117, 
                           ZN => n115);
   U161 : NAND2_X1 port map( A1 => n2371, A2 => n2407, ZN => n117);
   U162 : AOI221_X1 port map( B1 => DATA1(4), B2 => n2393, C1 => n2369, C2 => 
                           n2414, A => n2390, ZN => n116);
   U163 : INV_X1 port map( A => DATA1(4), ZN => n2414);
   U164 : OAI22_X1 port map( A1 => n111, A2 => n2415, B1 => n2442, B2 => n112, 
                           ZN => n110);
   U165 : NAND2_X1 port map( A1 => n2371, A2 => n2415, ZN => n112);
   U166 : INV_X1 port map( A => DATA1(5), ZN => n2415);
   U167 : AOI221_X1 port map( B1 => DATA2(5), B2 => n2393, C1 => n2369, C2 => 
                           n2442, A => n2390, ZN => n111);
   U168 : OAI22_X1 port map( A1 => n106_port, A2 => n2416, B1 => n2443, B2 => 
                           n107_port, ZN => n105_port);
   U169 : NAND2_X1 port map( A1 => n2371, A2 => n2416, ZN => n107_port);
   U170 : INV_X1 port map( A => DATA1(6), ZN => n2416);
   U171 : AOI221_X1 port map( B1 => DATA2(6), B2 => n2393, C1 => n2369, C2 => 
                           n2443, A => n2390, ZN => n106_port);
   U172 : OAI22_X1 port map( A1 => n101_port, A2 => n2417, B1 => n2444, B2 => 
                           n102_port, ZN => n100_port);
   U173 : NAND2_X1 port map( A1 => n2371, A2 => n2417, ZN => n102_port);
   U174 : INV_X1 port map( A => DATA1(7), ZN => n2417);
   U175 : AOI221_X1 port map( B1 => DATA2(7), B2 => n2393, C1 => n2368, C2 => 
                           n2444, A => n2390, ZN => n101_port);
   U176 : OAI22_X1 port map( A1 => n96_port, A2 => n2418, B1 => n2445, B2 => 
                           n97_port, ZN => n95_port);
   U177 : NAND2_X1 port map( A1 => n2370, A2 => n2418, ZN => n97_port);
   U178 : INV_X1 port map( A => DATA1(8), ZN => n2418);
   U179 : AOI221_X1 port map( B1 => DATA2(8), B2 => n2393, C1 => n2368, C2 => 
                           n2445, A => n2390, ZN => n96_port);
   U180 : OAI22_X1 port map( A1 => n86_port, A2 => n2419, B1 => n2446, B2 => 
                           n87_port, ZN => n85_port);
   U181 : NAND2_X1 port map( A1 => n2371, A2 => n2419, ZN => n87_port);
   U182 : INV_X1 port map( A => DATA1(9), ZN => n2419);
   U183 : AOI221_X1 port map( B1 => n2393, B2 => DATA2(9), C1 => n2368, C2 => 
                           n2446, A => n2390, ZN => n86_port);
   U184 : OAI22_X1 port map( A1 => n241, A2 => n2420, B1 => n2447, B2 => n242, 
                           ZN => n240);
   U185 : NAND2_X1 port map( A1 => n2371, A2 => n2420, ZN => n242);
   U186 : INV_X1 port map( A => DATA1(10), ZN => n2420);
   U187 : AOI221_X1 port map( B1 => DATA2(10), B2 => n2393, C1 => n2368, C2 => 
                           n2447, A => n2388, ZN => n241);
   U188 : OAI22_X1 port map( A1 => n236, A2 => n2421, B1 => n2448, B2 => n237, 
                           ZN => n235);
   U189 : NAND2_X1 port map( A1 => n2373, A2 => n2421, ZN => n237);
   U190 : INV_X1 port map( A => DATA1(11), ZN => n2421);
   U191 : AOI221_X1 port map( B1 => DATA2(11), B2 => n2395, C1 => n2368, C2 => 
                           n2448, A => n2388, ZN => n236);
   U192 : OAI22_X1 port map( A1 => n231, A2 => n2422, B1 => n2449, B2 => n232, 
                           ZN => n230);
   U193 : NAND2_X1 port map( A1 => n2373, A2 => n2422, ZN => n232);
   U194 : INV_X1 port map( A => DATA1(12), ZN => n2422);
   U195 : AOI221_X1 port map( B1 => DATA2(12), B2 => n2395, C1 => n2368, C2 => 
                           n2449, A => n2388, ZN => n231);
   U196 : OAI22_X1 port map( A1 => n226, A2 => n2450, B1 => n2423, B2 => n227, 
                           ZN => n225);
   U197 : NAND2_X1 port map( A1 => n2373, A2 => n2450, ZN => n227);
   U198 : INV_X1 port map( A => DATA2(13), ZN => n2450);
   U199 : AOI221_X1 port map( B1 => DATA1(13), B2 => n2395, C1 => n2368, C2 => 
                           n2423, A => n2388, ZN => n226);
   U200 : OAI22_X1 port map( A1 => n221, A2 => n2451, B1 => n2424, B2 => n222, 
                           ZN => n220);
   U201 : NAND2_X1 port map( A1 => n2373, A2 => n2451, ZN => n222);
   U202 : INV_X1 port map( A => DATA2(14), ZN => n2451);
   U203 : AOI221_X1 port map( B1 => DATA1(14), B2 => n2395, C1 => n2368, C2 => 
                           n2424, A => n2388, ZN => n221);
   U204 : OAI22_X1 port map( A1 => n216, A2 => n2452, B1 => n2425, B2 => n217, 
                           ZN => n215);
   U205 : NAND2_X1 port map( A1 => n2373, A2 => n2452, ZN => n217);
   U206 : INV_X1 port map( A => DATA2(15), ZN => n2452);
   U207 : AOI221_X1 port map( B1 => DATA1(15), B2 => n2395, C1 => n2368, C2 => 
                           n2425, A => n2388, ZN => n216);
   U208 : OAI22_X1 port map( A1 => n211, A2 => n2453, B1 => n2426, B2 => n212, 
                           ZN => n210);
   U209 : NAND2_X1 port map( A1 => n2373, A2 => n2453, ZN => n212);
   U210 : INV_X1 port map( A => DATA2(16), ZN => n2453);
   U211 : AOI221_X1 port map( B1 => DATA1(16), B2 => n2395, C1 => n2368, C2 => 
                           n2426, A => n2388, ZN => n211);
   U212 : OAI22_X1 port map( A1 => n206, A2 => n2454, B1 => n2427, B2 => n207, 
                           ZN => n205);
   U213 : NAND2_X1 port map( A1 => n2372, A2 => n2454, ZN => n207);
   U214 : INV_X1 port map( A => DATA2(17), ZN => n2454);
   U215 : AOI221_X1 port map( B1 => DATA1(17), B2 => n2395, C1 => n2369, C2 => 
                           n2427, A => n2388, ZN => n206);
   U216 : OAI22_X1 port map( A1 => n201, A2 => n2455, B1 => n2428, B2 => n202, 
                           ZN => n200);
   U217 : NAND2_X1 port map( A1 => n2372, A2 => n2455, ZN => n202);
   U218 : INV_X1 port map( A => DATA2(18), ZN => n2455);
   U219 : AOI221_X1 port map( B1 => DATA1(18), B2 => n2395, C1 => n2368, C2 => 
                           n2428, A => n2388, ZN => n201);
   U220 : OAI22_X1 port map( A1 => n196, A2 => n2456, B1 => n2429, B2 => n197, 
                           ZN => n195);
   U221 : NAND2_X1 port map( A1 => n2372, A2 => n2456, ZN => n197);
   U222 : INV_X1 port map( A => DATA2(19), ZN => n2456);
   U223 : AOI221_X1 port map( B1 => DATA1(19), B2 => n2394, C1 => n2369, C2 => 
                           n2429, A => n2388, ZN => n196);
   U224 : OAI22_X1 port map( A1 => n186, A2 => n2457, B1 => n2430, B2 => n187, 
                           ZN => n185);
   U225 : NAND2_X1 port map( A1 => n2372, A2 => n2457, ZN => n187);
   U226 : INV_X1 port map( A => DATA2(20), ZN => n2457);
   U227 : AOI221_X1 port map( B1 => DATA1(20), B2 => n2394, C1 => n2369, C2 => 
                           n2430, A => n2389, ZN => n186);
   U228 : OAI22_X1 port map( A1 => n181, A2 => n2431, B1 => n2458, B2 => n182, 
                           ZN => n180);
   U229 : NAND2_X1 port map( A1 => n2372, A2 => n2431, ZN => n182);
   U230 : INV_X1 port map( A => DATA1(21), ZN => n2431);
   U231 : AOI221_X1 port map( B1 => DATA2(21), B2 => n2394, C1 => n2369, C2 => 
                           n2458, A => n2389, ZN => n181);
   U232 : OAI22_X1 port map( A1 => n176, A2 => n2459, B1 => n2432, B2 => n177, 
                           ZN => n175);
   U233 : NAND2_X1 port map( A1 => n2372, A2 => n2459, ZN => n177);
   U234 : INV_X1 port map( A => DATA2(22), ZN => n2459);
   U235 : AOI221_X1 port map( B1 => DATA1(22), B2 => n2394, C1 => n2370, C2 => 
                           n2432, A => n2389, ZN => n176);
   U236 : OAI22_X1 port map( A1 => n171_port, A2 => n2433, B1 => n2460, B2 => 
                           n172_port, ZN => n170_port);
   U237 : NAND2_X1 port map( A1 => n2372, A2 => n2433, ZN => n172_port);
   U238 : INV_X1 port map( A => DATA1(23), ZN => n2433);
   U239 : AOI221_X1 port map( B1 => DATA2(23), B2 => n2394, C1 => n2369, C2 => 
                           n2460, A => n2389, ZN => n171_port);
   U240 : OAI22_X1 port map( A1 => n166_port, A2 => n2461, B1 => n2434, B2 => 
                           n167_port, ZN => n165_port);
   U241 : NAND2_X1 port map( A1 => n2372, A2 => n2461, ZN => n167_port);
   U242 : INV_X1 port map( A => DATA2(24), ZN => n2461);
   U243 : AOI221_X1 port map( B1 => DATA1(24), B2 => n2394, C1 => n2370, C2 => 
                           n2434, A => n2389, ZN => n166_port);
   U244 : OAI22_X1 port map( A1 => n161_port, A2 => n2435, B1 => n2462, B2 => 
                           n162_port, ZN => n160_port);
   U245 : NAND2_X1 port map( A1 => n2372, A2 => n2435, ZN => n162_port);
   U246 : INV_X1 port map( A => DATA1(25), ZN => n2435);
   U247 : AOI221_X1 port map( B1 => DATA2(25), B2 => n2394, C1 => n2370, C2 => 
                           n2462, A => n2389, ZN => n161_port);
   U248 : OAI22_X1 port map( A1 => n156_port, A2 => n2436, B1 => n2463, B2 => 
                           n157_port, ZN => n155_port);
   U249 : NAND2_X1 port map( A1 => n2372, A2 => n2436, ZN => n157_port);
   U250 : INV_X1 port map( A => DATA1(26), ZN => n2436);
   U251 : AOI221_X1 port map( B1 => DATA2(26), B2 => n2394, C1 => n2369, C2 => 
                           n2463, A => n2389, ZN => n156_port);
   U252 : OAI22_X1 port map( A1 => n151_port, A2 => n2437, B1 => n2464, B2 => 
                           n152_port, ZN => n150_port);
   U253 : NAND2_X1 port map( A1 => n2372, A2 => n2437, ZN => n152_port);
   U254 : INV_X1 port map( A => DATA1(27), ZN => n2437);
   U255 : AOI221_X1 port map( B1 => DATA2(27), B2 => n2394, C1 => n2370, C2 => 
                           n2464, A => n2389, ZN => n151_port);
   U256 : OAI22_X1 port map( A1 => n146_port, A2 => n2465, B1 => n2438, B2 => 
                           n147_port, ZN => n145_port);
   U257 : NAND2_X1 port map( A1 => n2371, A2 => n2465, ZN => n147_port);
   U258 : INV_X1 port map( A => DATA2(28), ZN => n2465);
   U259 : AOI221_X1 port map( B1 => DATA1(28), B2 => n2394, C1 => n2370, C2 => 
                           n2438, A => n2389, ZN => n146_port);
   U260 : OAI22_X1 port map( A1 => n141, A2 => n2439, B1 => n2466, B2 => 
                           n142_port, ZN => n140);
   U261 : NAND2_X1 port map( A1 => n2371, A2 => n2439, ZN => n142_port);
   U262 : INV_X1 port map( A => DATA1(29), ZN => n2439);
   U263 : AOI221_X1 port map( B1 => DATA2(29), B2 => n2393, C1 => n2370, C2 => 
                           n2466, A => n2389, ZN => n141);
   U264 : OAI22_X1 port map( A1 => n131, A2 => n2467, B1 => n2440, B2 => n132, 
                           ZN => n130);
   U265 : NAND2_X1 port map( A1 => n2371, A2 => n2467, ZN => n132);
   U266 : INV_X1 port map( A => DATA2(30), ZN => n2467);
   U267 : AOI221_X1 port map( B1 => DATA1(30), B2 => n2394, C1 => n2370, C2 => 
                           n2440, A => n2389, ZN => n131);
   U268 : OAI22_X1 port map( A1 => n126, A2 => n2441, B1 => n2468, B2 => n127, 
                           ZN => n125);
   U269 : NAND2_X1 port map( A1 => n2371, A2 => n2441, ZN => n127);
   U270 : INV_X1 port map( A => DATA1(31), ZN => n2441);
   U271 : AOI221_X1 port map( B1 => DATA2(31), B2 => n2393, C1 => n2369, C2 => 
                           n2468, A => n2390, ZN => n126);
   U272 : NOR2_X1 port map( A1 => FUNC(1), A2 => FUNC(0), ZN => n262);
   U273 : INV_X1 port map( A => FUNC(2), ZN => n2472);
   U274 : OAI21_X1 port map( B1 => n251, B2 => n252, A => FUNC(3), ZN => n250);
   U275 : NAND4_X1 port map( A1 => n253, A2 => n254, A3 => n255, A4 => n256, ZN
                           => n252);
   U276 : NAND4_X1 port map( A1 => n257, A2 => n258, A3 => n259, A4 => n260, ZN
                           => n251);
   U277 : NOR3_X1 port map( A1 => tmp_sub_0_port, A2 => tmp_sub_11_port, A3 => 
                           tmp_sub_10_port, ZN => n253);
   U278 : INV_X1 port map( A => FUNC(1), ZN => n2471);
   U279 : INV_X1 port map( A => FUNC(3), ZN => n2473);
   U280 : NOR4_X1 port map( A1 => n2472, A2 => n2471, A3 => FUNC(3), A4 => 
                           FUNC(0), ZN => n84_port);
   U281 : NOR4_X1 port map( A1 => n2472, A2 => n2473, A3 => n2471, A4 => 
                           FUNC(0), ZN => n83_port);
   U282 : NAND2_X1 port map( A1 => n123, A2 => n124, ZN => OUTALU(31));
   U283 : AOI221_X1 port map( B1 => N333, B2 => n2401, C1 => N301, C2 => n2396,
                           A => n125, ZN => n124);
   U284 : AOI222_X1 port map( A1 => N109, A2 => n2387, B1 => N173, B2 => n2383,
                           C1 => tmp_sub_31_port, C2 => n2379, ZN => n123);
   U285 : INV_X1 port map( A => DATA2(5), ZN => n2442);
   U286 : INV_X1 port map( A => DATA2(6), ZN => n2443);
   U287 : INV_X1 port map( A => DATA2(7), ZN => n2444);
   U288 : INV_X1 port map( A => DATA2(8), ZN => n2445);
   U289 : INV_X1 port map( A => DATA2(9), ZN => n2446);
   U290 : INV_X1 port map( A => DATA2(10), ZN => n2447);
   U291 : INV_X1 port map( A => DATA2(11), ZN => n2448);
   U292 : INV_X1 port map( A => DATA2(12), ZN => n2449);
   U296 : INV_X1 port map( A => DATA1(13), ZN => n2423);
   U297 : INV_X1 port map( A => DATA1(14), ZN => n2424);
   U298 : INV_X1 port map( A => DATA1(15), ZN => n2425);
   U299 : INV_X1 port map( A => DATA1(16), ZN => n2426);
   U300 : INV_X1 port map( A => DATA1(17), ZN => n2427);
   U301 : INV_X1 port map( A => DATA1(18), ZN => n2428);
   U302 : INV_X1 port map( A => DATA1(19), ZN => n2429);
   U303 : INV_X1 port map( A => DATA1(20), ZN => n2430);
   U304 : INV_X1 port map( A => DATA2(21), ZN => n2458);
   U305 : INV_X1 port map( A => DATA1(22), ZN => n2432);
   U306 : INV_X1 port map( A => DATA2(23), ZN => n2460);
   U307 : INV_X1 port map( A => DATA1(24), ZN => n2434);
   U308 : INV_X1 port map( A => DATA2(25), ZN => n2462);
   U309 : INV_X1 port map( A => DATA2(26), ZN => n2463);
   U310 : INV_X1 port map( A => DATA2(27), ZN => n2464);
   U311 : INV_X1 port map( A => DATA1(28), ZN => n2438);
   U312 : INV_X1 port map( A => DATA2(29), ZN => n2466);
   U313 : INV_X1 port map( A => DATA1(30), ZN => n2440);
   U314 : INV_X1 port map( A => DATA2(31), ZN => n2468);
   U315 : NOR2_X1 port map( A1 => n247, A2 => FUNC(3), ZN => n89_port);
   U316 : INV_X1 port map( A => n261, ZN => n2409);
   U317 : AOI221_X1 port map( B1 => n2410, B2 => n2370, C1 => n2393, C2 => 
                           DATA1(0), A => n2388, ZN => n261);
   U318 : INV_X1 port map( A => FUNC(0), ZN => n2470);
   U319 : AND3_X1 port map( A1 => FUNC(3), A2 => n262, A3 => FUNC(2), ZN => 
                           n88_port);
   U320 : AND3_X1 port map( A1 => n262, A2 => n2472, A3 => FUNC(3), ZN => 
                           n92_port);
   U321 : AND3_X1 port map( A1 => n262, A2 => n2473, A3 => FUNC(2), ZN => 
                           n91_port);
   U322 : INV_X1 port map( A => DATA1(0), ZN => n2410);
   U323 : INV_X1 port map( A => DATA2(2), ZN => n2405);
   U324 : INV_X1 port map( A => DATA2(4), ZN => n2407);
   U325 : INV_X1 port map( A => DATA2(1), ZN => n2404);
   U326 : INV_X1 port map( A => DATA2(3), ZN => n2406);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity adder_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  res : out std_logic_vector 
         (31 downto 0));

end adder_NBIT32;

architecture SYN_beh of adder_NBIT32 is

   component adder_NBIT32_DW01_add_0_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1066 : std_logic;

begin
   
   n1 <= '0';
   add_17 : adder_NBIT32_DW01_add_0_DW01_add_1 port map( A(31) => A(31), A(30) 
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => n1, SUM(31) => res(31),
                           SUM(30) => res(30), SUM(29) => res(29), SUM(28) => 
                           res(28), SUM(27) => res(27), SUM(26) => res(26), 
                           SUM(25) => res(25), SUM(24) => res(24), SUM(23) => 
                           res(23), SUM(22) => res(22), SUM(21) => res(21), 
                           SUM(20) => res(20), SUM(19) => res(19), SUM(18) => 
                           res(18), SUM(17) => res(17), SUM(16) => res(16), 
                           SUM(15) => res(15), SUM(14) => res(14), SUM(13) => 
                           res(13), SUM(12) => res(12), SUM(11) => res(11), 
                           SUM(10) => res(10), SUM(9) => res(9), SUM(8) => 
                           res(8), SUM(7) => res(7), SUM(6) => res(6), SUM(5) 
                           => res(5), SUM(4) => res(4), SUM(3) => res(3), 
                           SUM(2) => res(2), SUM(1) => res(1), SUM(0) => res(0)
                           , CO => n_1066);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity sign_extend_NBIT26_NBIT_F32 is

   port( A : in std_logic_vector (25 downto 0);  res : out std_logic_vector (31
         downto 0));

end sign_extend_NBIT26_NBIT_F32;

architecture SYN_beh of sign_extend_NBIT26_NBIT_F32 is

begin
   res <= ( A(25), A(25), A(25), A(25), A(25), A(25), A(25), A(24), A(23), 
      A(22), A(21), A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), 
      A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1)
      , A(0) );

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity AND2 is

   port( a, b : in std_logic;  y : out std_logic);

end AND2;

architecture SYN_BEHAVIORAL of AND2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IV is

   port( A : in std_logic;  Y : out std_logic);

end IV;

architecture SYN_BEHAVIORAL of IV is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity sign_extend_NBIT16_NBIT_F32 is

   port( A : in std_logic_vector (15 downto 0);  res : out std_logic_vector (31
         downto 0));

end sign_extend_NBIT16_NBIT_F32;

architecture SYN_beh of sign_extend_NBIT16_NBIT_F32 is

begin
   res <= ( A(15), A(15), A(15), A(15), A(15), A(15), A(15), A(15), A(15), 
      A(15), A(15), A(15), A(15), A(15), A(15), A(15), A(15), A(14), A(13), 
      A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1)
      , A(0) );

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity reg_file_NBIT32_NREG32_NADDR5 is

   port( clk, rst, wr_en : in std_logic;  add_rd1, add_rd2 : in 
         std_logic_vector (4 downto 0);  add_wr, datain : in std_logic_vector 
         (31 downto 0);  out2, out1 : out std_logic_vector (31 downto 0));

end reg_file_NBIT32_NREG32_NADDR5;

architecture SYN_beh of reg_file_NBIT32_NREG32_NADDR5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal regs_5_31_port, regs_5_30_port, regs_5_29_port, regs_5_28_port, 
      regs_5_27_port, regs_5_26_port, regs_5_25_port, regs_5_24_port, 
      regs_5_23_port, regs_5_22_port, regs_5_21_port, regs_5_20_port, 
      regs_5_19_port, regs_5_18_port, regs_5_17_port, regs_5_16_port, 
      regs_5_15_port, regs_5_14_port, regs_5_13_port, regs_5_12_port, 
      regs_5_11_port, regs_5_10_port, regs_5_9_port, regs_5_8_port, 
      regs_5_7_port, regs_5_6_port, regs_5_5_port, regs_5_4_port, regs_5_3_port
      , regs_5_2_port, regs_5_1_port, regs_5_0_port, regs_7_31_port, 
      regs_7_30_port, regs_7_29_port, regs_7_28_port, regs_7_27_port, 
      regs_7_26_port, regs_7_25_port, regs_7_24_port, regs_7_23_port, 
      regs_7_22_port, regs_7_21_port, regs_7_20_port, regs_7_19_port, 
      regs_7_18_port, regs_7_17_port, regs_7_16_port, regs_7_15_port, 
      regs_7_14_port, regs_7_13_port, regs_7_12_port, regs_7_11_port, 
      regs_7_10_port, regs_7_9_port, regs_7_8_port, regs_7_7_port, 
      regs_7_6_port, regs_7_5_port, regs_7_4_port, regs_7_3_port, regs_7_2_port
      , regs_7_1_port, regs_7_0_port, regs_13_31_port, regs_13_30_port, 
      regs_13_29_port, regs_13_28_port, regs_13_27_port, regs_13_26_port, 
      regs_13_25_port, regs_13_24_port, regs_13_23_port, regs_13_22_port, 
      regs_13_21_port, regs_13_20_port, regs_13_19_port, regs_13_18_port, 
      regs_13_17_port, regs_13_16_port, regs_13_15_port, regs_13_14_port, 
      regs_13_13_port, regs_13_12_port, regs_13_11_port, regs_13_10_port, 
      regs_13_9_port, regs_13_8_port, regs_13_7_port, regs_13_6_port, 
      regs_13_5_port, regs_13_4_port, regs_13_3_port, regs_13_2_port, 
      regs_13_1_port, regs_13_0_port, regs_15_31_port, regs_15_30_port, 
      regs_15_29_port, regs_15_28_port, regs_15_27_port, regs_15_26_port, 
      regs_15_25_port, regs_15_24_port, regs_15_23_port, regs_15_22_port, 
      regs_15_21_port, regs_15_20_port, regs_15_19_port, regs_15_18_port, 
      regs_15_17_port, regs_15_16_port, regs_15_15_port, regs_15_14_port, 
      regs_15_13_port, regs_15_12_port, regs_15_11_port, regs_15_10_port, 
      regs_15_9_port, regs_15_8_port, regs_15_7_port, regs_15_6_port, 
      regs_15_5_port, regs_15_4_port, regs_15_3_port, regs_15_2_port, 
      regs_15_1_port, regs_15_0_port, regs_18_31_port, regs_18_30_port, 
      regs_18_29_port, regs_18_28_port, regs_18_27_port, regs_18_26_port, 
      regs_18_25_port, regs_18_24_port, regs_18_23_port, regs_18_22_port, 
      regs_18_21_port, regs_18_20_port, regs_18_19_port, regs_18_18_port, 
      regs_18_17_port, regs_18_16_port, regs_18_15_port, regs_18_14_port, 
      regs_18_13_port, regs_18_12_port, regs_18_11_port, regs_18_10_port, 
      regs_18_9_port, regs_18_8_port, regs_18_7_port, regs_18_6_port, 
      regs_18_5_port, regs_18_4_port, regs_18_3_port, regs_18_2_port, 
      regs_18_1_port, regs_18_0_port, regs_nxt_0_31_port, regs_nxt_0_30_port, 
      regs_nxt_0_29_port, regs_nxt_0_28_port, regs_nxt_0_27_port, 
      regs_nxt_0_26_port, regs_nxt_0_25_port, regs_nxt_0_24_port, 
      regs_nxt_0_23_port, regs_nxt_0_22_port, regs_nxt_0_21_port, 
      regs_nxt_0_20_port, regs_nxt_0_19_port, regs_nxt_0_18_port, 
      regs_nxt_0_17_port, regs_nxt_0_16_port, regs_nxt_0_15_port, 
      regs_nxt_0_14_port, regs_nxt_0_13_port, regs_nxt_0_12_port, 
      regs_nxt_0_11_port, regs_nxt_0_10_port, regs_nxt_0_9_port, 
      regs_nxt_0_8_port, regs_nxt_0_7_port, regs_nxt_0_6_port, 
      regs_nxt_0_5_port, regs_nxt_0_4_port, regs_nxt_0_3_port, 
      regs_nxt_0_2_port, regs_nxt_0_1_port, regs_nxt_0_0_port, 
      regs_nxt_1_31_port, regs_nxt_1_30_port, regs_nxt_1_29_port, 
      regs_nxt_1_28_port, regs_nxt_1_27_port, regs_nxt_1_26_port, 
      regs_nxt_1_25_port, regs_nxt_1_24_port, regs_nxt_1_23_port, 
      regs_nxt_1_22_port, regs_nxt_1_21_port, regs_nxt_1_20_port, 
      regs_nxt_1_19_port, regs_nxt_1_18_port, regs_nxt_1_17_port, 
      regs_nxt_1_16_port, regs_nxt_1_15_port, regs_nxt_1_14_port, 
      regs_nxt_1_13_port, regs_nxt_1_12_port, regs_nxt_1_11_port, 
      regs_nxt_1_10_port, regs_nxt_1_9_port, regs_nxt_1_8_port, 
      regs_nxt_1_7_port, regs_nxt_1_6_port, regs_nxt_1_5_port, 
      regs_nxt_1_4_port, regs_nxt_1_3_port, regs_nxt_1_2_port, 
      regs_nxt_1_1_port, regs_nxt_1_0_port, regs_nxt_2_31_port, 
      regs_nxt_2_30_port, regs_nxt_2_29_port, regs_nxt_2_28_port, 
      regs_nxt_2_27_port, regs_nxt_2_26_port, regs_nxt_2_25_port, 
      regs_nxt_2_24_port, regs_nxt_2_23_port, regs_nxt_2_22_port, 
      regs_nxt_2_21_port, regs_nxt_2_20_port, regs_nxt_2_19_port, 
      regs_nxt_2_18_port, regs_nxt_2_17_port, regs_nxt_2_16_port, 
      regs_nxt_2_15_port, regs_nxt_2_14_port, regs_nxt_2_13_port, 
      regs_nxt_2_12_port, regs_nxt_2_11_port, regs_nxt_2_10_port, 
      regs_nxt_2_9_port, regs_nxt_2_8_port, regs_nxt_2_7_port, 
      regs_nxt_2_6_port, regs_nxt_2_5_port, regs_nxt_2_4_port, 
      regs_nxt_2_3_port, regs_nxt_2_2_port, regs_nxt_2_1_port, 
      regs_nxt_2_0_port, regs_nxt_3_31_port, regs_nxt_3_30_port, 
      regs_nxt_3_29_port, regs_nxt_3_28_port, regs_nxt_3_27_port, 
      regs_nxt_3_26_port, regs_nxt_3_25_port, regs_nxt_3_24_port, 
      regs_nxt_3_23_port, regs_nxt_3_22_port, regs_nxt_3_21_port, 
      regs_nxt_3_20_port, regs_nxt_3_19_port, regs_nxt_3_18_port, 
      regs_nxt_3_17_port, regs_nxt_3_16_port, regs_nxt_3_15_port, 
      regs_nxt_3_14_port, regs_nxt_3_13_port, regs_nxt_3_12_port, 
      regs_nxt_3_11_port, regs_nxt_3_10_port, regs_nxt_3_9_port, 
      regs_nxt_3_8_port, regs_nxt_3_7_port, regs_nxt_3_6_port, 
      regs_nxt_3_5_port, regs_nxt_3_4_port, regs_nxt_3_3_port, 
      regs_nxt_3_2_port, regs_nxt_3_1_port, regs_nxt_3_0_port, 
      regs_nxt_4_31_port, regs_nxt_4_30_port, regs_nxt_4_29_port, 
      regs_nxt_4_28_port, regs_nxt_4_27_port, regs_nxt_4_26_port, 
      regs_nxt_4_25_port, regs_nxt_4_24_port, regs_nxt_4_23_port, 
      regs_nxt_4_22_port, regs_nxt_4_21_port, regs_nxt_4_20_port, 
      regs_nxt_4_19_port, regs_nxt_4_18_port, regs_nxt_4_17_port, 
      regs_nxt_4_16_port, regs_nxt_4_15_port, regs_nxt_4_14_port, 
      regs_nxt_4_13_port, regs_nxt_4_12_port, regs_nxt_4_11_port, 
      regs_nxt_4_10_port, regs_nxt_4_9_port, regs_nxt_4_8_port, 
      regs_nxt_4_7_port, regs_nxt_4_6_port, regs_nxt_4_5_port, 
      regs_nxt_4_4_port, regs_nxt_4_3_port, regs_nxt_4_2_port, 
      regs_nxt_4_1_port, regs_nxt_4_0_port, regs_nxt_5_31_port, 
      regs_nxt_5_30_port, regs_nxt_5_29_port, regs_nxt_5_28_port, 
      regs_nxt_5_27_port, regs_nxt_5_26_port, regs_nxt_5_25_port, 
      regs_nxt_5_24_port, regs_nxt_5_23_port, regs_nxt_5_22_port, 
      regs_nxt_5_21_port, regs_nxt_5_20_port, regs_nxt_5_19_port, 
      regs_nxt_5_18_port, regs_nxt_5_17_port, regs_nxt_5_16_port, 
      regs_nxt_5_15_port, regs_nxt_5_14_port, regs_nxt_5_13_port, 
      regs_nxt_5_12_port, regs_nxt_5_11_port, regs_nxt_5_10_port, 
      regs_nxt_5_9_port, regs_nxt_5_8_port, regs_nxt_5_7_port, 
      regs_nxt_5_6_port, regs_nxt_5_5_port, regs_nxt_5_4_port, 
      regs_nxt_5_3_port, regs_nxt_5_2_port, regs_nxt_5_1_port, 
      regs_nxt_5_0_port, regs_nxt_6_31_port, regs_nxt_6_30_port, 
      regs_nxt_6_29_port, regs_nxt_6_28_port, regs_nxt_6_27_port, 
      regs_nxt_6_26_port, regs_nxt_6_25_port, regs_nxt_6_24_port, 
      regs_nxt_6_23_port, regs_nxt_6_22_port, regs_nxt_6_21_port, 
      regs_nxt_6_20_port, regs_nxt_6_19_port, regs_nxt_6_18_port, 
      regs_nxt_6_17_port, regs_nxt_6_16_port, regs_nxt_6_15_port, 
      regs_nxt_6_14_port, regs_nxt_6_13_port, regs_nxt_6_12_port, 
      regs_nxt_6_11_port, regs_nxt_6_10_port, regs_nxt_6_9_port, 
      regs_nxt_6_8_port, regs_nxt_6_7_port, regs_nxt_6_6_port, 
      regs_nxt_6_5_port, regs_nxt_6_4_port, regs_nxt_6_3_port, 
      regs_nxt_6_2_port, regs_nxt_6_1_port, regs_nxt_6_0_port, 
      regs_nxt_7_31_port, regs_nxt_7_30_port, regs_nxt_7_29_port, 
      regs_nxt_7_28_port, regs_nxt_7_27_port, regs_nxt_7_26_port, 
      regs_nxt_7_25_port, regs_nxt_7_24_port, regs_nxt_7_23_port, 
      regs_nxt_7_22_port, regs_nxt_7_21_port, regs_nxt_7_20_port, 
      regs_nxt_7_19_port, regs_nxt_7_18_port, regs_nxt_7_17_port, 
      regs_nxt_7_16_port, regs_nxt_7_15_port, regs_nxt_7_14_port, 
      regs_nxt_7_13_port, regs_nxt_7_12_port, regs_nxt_7_11_port, 
      regs_nxt_7_10_port, regs_nxt_7_9_port, regs_nxt_7_8_port, 
      regs_nxt_7_7_port, regs_nxt_7_6_port, regs_nxt_7_5_port, 
      regs_nxt_7_4_port, regs_nxt_7_3_port, regs_nxt_7_2_port, 
      regs_nxt_7_1_port, regs_nxt_7_0_port, regs_nxt_8_31_port, 
      regs_nxt_8_30_port, regs_nxt_8_29_port, regs_nxt_8_28_port, 
      regs_nxt_8_27_port, regs_nxt_8_26_port, regs_nxt_8_25_port, 
      regs_nxt_8_24_port, regs_nxt_8_23_port, regs_nxt_8_22_port, 
      regs_nxt_8_21_port, regs_nxt_8_20_port, regs_nxt_8_19_port, 
      regs_nxt_8_18_port, regs_nxt_8_17_port, regs_nxt_8_16_port, 
      regs_nxt_8_15_port, regs_nxt_8_14_port, regs_nxt_8_13_port, 
      regs_nxt_8_12_port, regs_nxt_8_11_port, regs_nxt_8_10_port, 
      regs_nxt_8_9_port, regs_nxt_8_8_port, regs_nxt_8_7_port, 
      regs_nxt_8_6_port, regs_nxt_8_5_port, regs_nxt_8_4_port, 
      regs_nxt_8_3_port, regs_nxt_8_2_port, regs_nxt_8_1_port, 
      regs_nxt_8_0_port, regs_nxt_9_31_port, regs_nxt_9_30_port, 
      regs_nxt_9_29_port, regs_nxt_9_28_port, regs_nxt_9_27_port, 
      regs_nxt_9_26_port, regs_nxt_9_25_port, regs_nxt_9_24_port, 
      regs_nxt_9_23_port, regs_nxt_9_22_port, regs_nxt_9_21_port, 
      regs_nxt_9_20_port, regs_nxt_9_19_port, regs_nxt_9_18_port, 
      regs_nxt_9_17_port, regs_nxt_9_16_port, regs_nxt_9_15_port, 
      regs_nxt_9_14_port, regs_nxt_9_13_port, regs_nxt_9_12_port, 
      regs_nxt_9_11_port, regs_nxt_9_10_port, regs_nxt_9_9_port, 
      regs_nxt_9_8_port, regs_nxt_9_7_port, regs_nxt_9_6_port, 
      regs_nxt_9_5_port, regs_nxt_9_4_port, regs_nxt_9_3_port, 
      regs_nxt_9_2_port, regs_nxt_9_1_port, regs_nxt_9_0_port, 
      regs_nxt_10_31_port, regs_nxt_10_30_port, regs_nxt_10_29_port, 
      regs_nxt_10_28_port, regs_nxt_10_27_port, regs_nxt_10_26_port, 
      regs_nxt_10_25_port, regs_nxt_10_24_port, regs_nxt_10_23_port, 
      regs_nxt_10_22_port, regs_nxt_10_21_port, regs_nxt_10_20_port, 
      regs_nxt_10_19_port, regs_nxt_10_18_port, regs_nxt_10_17_port, 
      regs_nxt_10_16_port, regs_nxt_10_15_port, regs_nxt_10_14_port, 
      regs_nxt_10_13_port, regs_nxt_10_12_port, regs_nxt_10_11_port, 
      regs_nxt_10_10_port, regs_nxt_10_9_port, regs_nxt_10_8_port, 
      regs_nxt_10_7_port, regs_nxt_10_6_port, regs_nxt_10_5_port, 
      regs_nxt_10_4_port, regs_nxt_10_3_port, regs_nxt_10_2_port, 
      regs_nxt_10_1_port, regs_nxt_10_0_port, regs_nxt_11_31_port, 
      regs_nxt_11_30_port, regs_nxt_11_29_port, regs_nxt_11_28_port, 
      regs_nxt_11_27_port, regs_nxt_11_26_port, regs_nxt_11_25_port, 
      regs_nxt_11_24_port, regs_nxt_11_23_port, regs_nxt_11_22_port, 
      regs_nxt_11_21_port, regs_nxt_11_20_port, regs_nxt_11_19_port, 
      regs_nxt_11_18_port, regs_nxt_11_17_port, regs_nxt_11_16_port, 
      regs_nxt_11_15_port, regs_nxt_11_14_port, regs_nxt_11_13_port, 
      regs_nxt_11_12_port, regs_nxt_11_11_port, regs_nxt_11_10_port, 
      regs_nxt_11_9_port, regs_nxt_11_8_port, regs_nxt_11_7_port, 
      regs_nxt_11_6_port, regs_nxt_11_5_port, regs_nxt_11_4_port, 
      regs_nxt_11_3_port, regs_nxt_11_2_port, regs_nxt_11_1_port, 
      regs_nxt_11_0_port, regs_nxt_12_31_port, regs_nxt_12_30_port, 
      regs_nxt_12_29_port, regs_nxt_12_28_port, regs_nxt_12_27_port, 
      regs_nxt_12_26_port, regs_nxt_12_25_port, regs_nxt_12_24_port, 
      regs_nxt_12_23_port, regs_nxt_12_22_port, regs_nxt_12_21_port, 
      regs_nxt_12_20_port, regs_nxt_12_19_port, regs_nxt_12_18_port, 
      regs_nxt_12_17_port, regs_nxt_12_16_port, regs_nxt_12_15_port, 
      regs_nxt_12_14_port, regs_nxt_12_13_port, regs_nxt_12_12_port, 
      regs_nxt_12_11_port, regs_nxt_12_10_port, regs_nxt_12_9_port, 
      regs_nxt_12_8_port, regs_nxt_12_7_port, regs_nxt_12_6_port, 
      regs_nxt_12_5_port, regs_nxt_12_4_port, regs_nxt_12_3_port, 
      regs_nxt_12_2_port, regs_nxt_12_1_port, regs_nxt_12_0_port, 
      regs_nxt_13_31_port, regs_nxt_13_30_port, regs_nxt_13_29_port, 
      regs_nxt_13_28_port, regs_nxt_13_27_port, regs_nxt_13_26_port, 
      regs_nxt_13_25_port, regs_nxt_13_24_port, regs_nxt_13_23_port, 
      regs_nxt_13_22_port, regs_nxt_13_21_port, regs_nxt_13_20_port, 
      regs_nxt_13_19_port, regs_nxt_13_18_port, regs_nxt_13_17_port, 
      regs_nxt_13_16_port, regs_nxt_13_15_port, regs_nxt_13_14_port, 
      regs_nxt_13_13_port, regs_nxt_13_12_port, regs_nxt_13_11_port, 
      regs_nxt_13_10_port, regs_nxt_13_9_port, regs_nxt_13_8_port, 
      regs_nxt_13_7_port, regs_nxt_13_6_port, regs_nxt_13_5_port, 
      regs_nxt_13_4_port, regs_nxt_13_3_port, regs_nxt_13_2_port, 
      regs_nxt_13_1_port, regs_nxt_13_0_port, regs_nxt_14_31_port, 
      regs_nxt_14_30_port, regs_nxt_14_29_port, regs_nxt_14_28_port, 
      regs_nxt_14_27_port, regs_nxt_14_26_port, regs_nxt_14_25_port, 
      regs_nxt_14_24_port, regs_nxt_14_23_port, regs_nxt_14_22_port, 
      regs_nxt_14_21_port, regs_nxt_14_20_port, regs_nxt_14_19_port, 
      regs_nxt_14_18_port, regs_nxt_14_17_port, regs_nxt_14_16_port, 
      regs_nxt_14_15_port, regs_nxt_14_14_port, regs_nxt_14_13_port, 
      regs_nxt_14_12_port, regs_nxt_14_11_port, regs_nxt_14_10_port, 
      regs_nxt_14_9_port, regs_nxt_14_8_port, regs_nxt_14_7_port, 
      regs_nxt_14_6_port, regs_nxt_14_5_port, regs_nxt_14_4_port, 
      regs_nxt_14_3_port, regs_nxt_14_2_port, regs_nxt_14_1_port, 
      regs_nxt_14_0_port, regs_nxt_15_31_port, regs_nxt_15_30_port, 
      regs_nxt_15_29_port, regs_nxt_15_28_port, regs_nxt_15_27_port, 
      regs_nxt_15_26_port, regs_nxt_15_25_port, regs_nxt_15_24_port, 
      regs_nxt_15_23_port, regs_nxt_15_22_port, regs_nxt_15_21_port, 
      regs_nxt_15_20_port, regs_nxt_15_19_port, regs_nxt_15_18_port, 
      regs_nxt_15_17_port, regs_nxt_15_16_port, regs_nxt_15_15_port, 
      regs_nxt_15_14_port, regs_nxt_15_13_port, regs_nxt_15_12_port, 
      regs_nxt_15_11_port, regs_nxt_15_10_port, regs_nxt_15_9_port, 
      regs_nxt_15_8_port, regs_nxt_15_7_port, regs_nxt_15_6_port, 
      regs_nxt_15_5_port, regs_nxt_15_4_port, regs_nxt_15_3_port, 
      regs_nxt_15_2_port, regs_nxt_15_1_port, regs_nxt_15_0_port, 
      regs_nxt_16_31_port, regs_nxt_16_30_port, regs_nxt_16_29_port, 
      regs_nxt_16_28_port, regs_nxt_16_27_port, regs_nxt_16_26_port, 
      regs_nxt_16_25_port, regs_nxt_16_24_port, regs_nxt_16_23_port, 
      regs_nxt_16_22_port, regs_nxt_16_21_port, regs_nxt_16_20_port, 
      regs_nxt_16_19_port, regs_nxt_16_18_port, regs_nxt_16_17_port, 
      regs_nxt_16_16_port, regs_nxt_16_15_port, regs_nxt_16_14_port, 
      regs_nxt_16_13_port, regs_nxt_16_12_port, regs_nxt_16_11_port, 
      regs_nxt_16_10_port, regs_nxt_16_9_port, regs_nxt_16_8_port, 
      regs_nxt_16_7_port, regs_nxt_16_6_port, regs_nxt_16_5_port, 
      regs_nxt_16_4_port, regs_nxt_16_3_port, regs_nxt_16_2_port, 
      regs_nxt_16_1_port, regs_nxt_16_0_port, regs_nxt_17_31_port, 
      regs_nxt_17_30_port, regs_nxt_17_29_port, regs_nxt_17_28_port, 
      regs_nxt_17_27_port, regs_nxt_17_26_port, regs_nxt_17_25_port, 
      regs_nxt_17_24_port, regs_nxt_17_23_port, regs_nxt_17_22_port, 
      regs_nxt_17_21_port, regs_nxt_17_20_port, regs_nxt_17_19_port, 
      regs_nxt_17_18_port, regs_nxt_17_17_port, regs_nxt_17_16_port, 
      regs_nxt_17_15_port, regs_nxt_17_14_port, regs_nxt_17_13_port, 
      regs_nxt_17_12_port, regs_nxt_17_11_port, regs_nxt_17_10_port, 
      regs_nxt_17_9_port, regs_nxt_17_8_port, regs_nxt_17_7_port, 
      regs_nxt_17_6_port, regs_nxt_17_5_port, regs_nxt_17_4_port, 
      regs_nxt_17_3_port, regs_nxt_17_2_port, regs_nxt_17_1_port, 
      regs_nxt_17_0_port, regs_nxt_18_31_port, regs_nxt_18_30_port, 
      regs_nxt_18_29_port, regs_nxt_18_28_port, regs_nxt_18_27_port, 
      regs_nxt_18_26_port, regs_nxt_18_25_port, regs_nxt_18_24_port, 
      regs_nxt_18_23_port, regs_nxt_18_22_port, regs_nxt_18_21_port, 
      regs_nxt_18_20_port, regs_nxt_18_19_port, regs_nxt_18_18_port, 
      regs_nxt_18_17_port, regs_nxt_18_16_port, regs_nxt_18_15_port, 
      regs_nxt_18_14_port, regs_nxt_18_13_port, regs_nxt_18_12_port, 
      regs_nxt_18_11_port, regs_nxt_18_10_port, regs_nxt_18_9_port, 
      regs_nxt_18_8_port, regs_nxt_18_7_port, regs_nxt_18_6_port, 
      regs_nxt_18_5_port, regs_nxt_18_4_port, regs_nxt_18_3_port, 
      regs_nxt_18_2_port, regs_nxt_18_1_port, regs_nxt_18_0_port, 
      regs_nxt_19_31_port, regs_nxt_19_30_port, regs_nxt_19_29_port, 
      regs_nxt_19_28_port, regs_nxt_19_27_port, regs_nxt_19_26_port, 
      regs_nxt_19_25_port, regs_nxt_19_24_port, regs_nxt_19_23_port, 
      regs_nxt_19_22_port, regs_nxt_19_21_port, regs_nxt_19_20_port, 
      regs_nxt_19_19_port, regs_nxt_19_18_port, regs_nxt_19_17_port, 
      regs_nxt_19_16_port, regs_nxt_19_15_port, regs_nxt_19_14_port, 
      regs_nxt_19_13_port, regs_nxt_19_12_port, regs_nxt_19_11_port, 
      regs_nxt_19_10_port, regs_nxt_19_9_port, regs_nxt_19_8_port, 
      regs_nxt_19_7_port, regs_nxt_19_6_port, regs_nxt_19_5_port, 
      regs_nxt_19_4_port, regs_nxt_19_3_port, regs_nxt_19_2_port, 
      regs_nxt_19_1_port, regs_nxt_19_0_port, regs_nxt_20_31_port, 
      regs_nxt_20_30_port, regs_nxt_20_29_port, regs_nxt_20_28_port, 
      regs_nxt_20_27_port, regs_nxt_20_26_port, regs_nxt_20_25_port, 
      regs_nxt_20_24_port, regs_nxt_20_23_port, regs_nxt_20_22_port, 
      regs_nxt_20_21_port, regs_nxt_20_20_port, regs_nxt_20_19_port, 
      regs_nxt_20_18_port, regs_nxt_20_17_port, regs_nxt_20_16_port, 
      regs_nxt_20_15_port, regs_nxt_20_14_port, regs_nxt_20_13_port, 
      regs_nxt_20_12_port, regs_nxt_20_11_port, regs_nxt_20_10_port, 
      regs_nxt_20_9_port, regs_nxt_20_8_port, regs_nxt_20_7_port, 
      regs_nxt_20_6_port, regs_nxt_20_5_port, regs_nxt_20_4_port, 
      regs_nxt_20_3_port, regs_nxt_20_2_port, regs_nxt_20_1_port, 
      regs_nxt_20_0_port, regs_nxt_21_31_port, regs_nxt_21_30_port, 
      regs_nxt_21_29_port, regs_nxt_21_28_port, regs_nxt_21_27_port, 
      regs_nxt_21_26_port, regs_nxt_21_25_port, regs_nxt_21_24_port, 
      regs_nxt_21_23_port, regs_nxt_21_22_port, regs_nxt_21_21_port, 
      regs_nxt_21_20_port, regs_nxt_21_19_port, regs_nxt_21_18_port, 
      regs_nxt_21_17_port, regs_nxt_21_16_port, regs_nxt_21_15_port, 
      regs_nxt_21_14_port, regs_nxt_21_13_port, regs_nxt_21_12_port, 
      regs_nxt_21_11_port, regs_nxt_21_10_port, regs_nxt_21_9_port, 
      regs_nxt_21_8_port, regs_nxt_21_7_port, regs_nxt_21_6_port, 
      regs_nxt_21_5_port, regs_nxt_21_4_port, regs_nxt_21_3_port, 
      regs_nxt_21_2_port, regs_nxt_21_1_port, regs_nxt_21_0_port, 
      regs_nxt_22_31_port, regs_nxt_22_30_port, regs_nxt_22_29_port, 
      regs_nxt_22_28_port, regs_nxt_22_27_port, regs_nxt_22_26_port, 
      regs_nxt_22_25_port, regs_nxt_22_24_port, regs_nxt_22_23_port, 
      regs_nxt_22_22_port, regs_nxt_22_21_port, regs_nxt_22_20_port, 
      regs_nxt_22_19_port, regs_nxt_22_18_port, regs_nxt_22_17_port, 
      regs_nxt_22_16_port, regs_nxt_22_15_port, regs_nxt_22_14_port, 
      regs_nxt_22_13_port, regs_nxt_22_12_port, regs_nxt_22_11_port, 
      regs_nxt_22_10_port, regs_nxt_22_9_port, regs_nxt_22_8_port, 
      regs_nxt_22_7_port, regs_nxt_22_6_port, regs_nxt_22_5_port, 
      regs_nxt_22_4_port, regs_nxt_22_3_port, regs_nxt_22_2_port, 
      regs_nxt_22_1_port, regs_nxt_22_0_port, regs_nxt_23_31_port, 
      regs_nxt_23_30_port, regs_nxt_23_29_port, regs_nxt_23_28_port, 
      regs_nxt_23_27_port, regs_nxt_23_26_port, regs_nxt_23_25_port, 
      regs_nxt_23_24_port, regs_nxt_23_23_port, regs_nxt_23_22_port, 
      regs_nxt_23_21_port, regs_nxt_23_20_port, regs_nxt_23_19_port, 
      regs_nxt_23_18_port, regs_nxt_23_17_port, regs_nxt_23_16_port, 
      regs_nxt_23_15_port, regs_nxt_23_14_port, regs_nxt_23_13_port, 
      regs_nxt_23_12_port, regs_nxt_23_11_port, regs_nxt_23_10_port, 
      regs_nxt_23_9_port, regs_nxt_23_8_port, regs_nxt_23_7_port, 
      regs_nxt_23_6_port, regs_nxt_23_5_port, regs_nxt_23_4_port, 
      regs_nxt_23_3_port, regs_nxt_23_2_port, regs_nxt_23_1_port, 
      regs_nxt_23_0_port, regs_nxt_24_31_port, regs_nxt_24_30_port, 
      regs_nxt_24_29_port, regs_nxt_24_28_port, regs_nxt_24_27_port, 
      regs_nxt_24_26_port, regs_nxt_24_25_port, regs_nxt_24_24_port, 
      regs_nxt_24_23_port, regs_nxt_24_22_port, regs_nxt_24_21_port, 
      regs_nxt_24_20_port, regs_nxt_24_19_port, regs_nxt_24_18_port, 
      regs_nxt_24_17_port, regs_nxt_24_16_port, regs_nxt_24_15_port, 
      regs_nxt_24_14_port, regs_nxt_24_13_port, regs_nxt_24_12_port, 
      regs_nxt_24_11_port, regs_nxt_24_10_port, regs_nxt_24_9_port, 
      regs_nxt_24_8_port, regs_nxt_24_7_port, regs_nxt_24_6_port, 
      regs_nxt_24_5_port, regs_nxt_24_4_port, regs_nxt_24_3_port, 
      regs_nxt_24_2_port, regs_nxt_24_1_port, regs_nxt_24_0_port, 
      regs_nxt_25_31_port, regs_nxt_25_30_port, regs_nxt_25_29_port, 
      regs_nxt_25_28_port, regs_nxt_25_27_port, regs_nxt_25_26_port, 
      regs_nxt_25_25_port, regs_nxt_25_24_port, regs_nxt_25_23_port, 
      regs_nxt_25_22_port, regs_nxt_25_21_port, regs_nxt_25_20_port, 
      regs_nxt_25_19_port, regs_nxt_25_18_port, regs_nxt_25_17_port, 
      regs_nxt_25_16_port, regs_nxt_25_15_port, regs_nxt_25_14_port, 
      regs_nxt_25_13_port, regs_nxt_25_12_port, regs_nxt_25_11_port, 
      regs_nxt_25_10_port, regs_nxt_25_9_port, regs_nxt_25_8_port, 
      regs_nxt_25_7_port, regs_nxt_25_6_port, regs_nxt_25_5_port, 
      regs_nxt_25_4_port, regs_nxt_25_3_port, regs_nxt_25_2_port, 
      regs_nxt_25_1_port, regs_nxt_25_0_port, regs_nxt_26_31_port, 
      regs_nxt_26_30_port, regs_nxt_26_29_port, regs_nxt_26_28_port, 
      regs_nxt_26_27_port, regs_nxt_26_26_port, regs_nxt_26_25_port, 
      regs_nxt_26_24_port, regs_nxt_26_23_port, regs_nxt_26_22_port, 
      regs_nxt_26_21_port, regs_nxt_26_20_port, regs_nxt_26_19_port, 
      regs_nxt_26_18_port, regs_nxt_26_17_port, regs_nxt_26_16_port, 
      regs_nxt_26_15_port, regs_nxt_26_14_port, regs_nxt_26_13_port, 
      regs_nxt_26_12_port, regs_nxt_26_11_port, regs_nxt_26_10_port, 
      regs_nxt_26_9_port, regs_nxt_26_8_port, regs_nxt_26_7_port, 
      regs_nxt_26_6_port, regs_nxt_26_5_port, regs_nxt_26_4_port, 
      regs_nxt_26_3_port, regs_nxt_26_2_port, regs_nxt_26_1_port, 
      regs_nxt_26_0_port, regs_nxt_27_31_port, regs_nxt_27_30_port, 
      regs_nxt_27_29_port, regs_nxt_27_28_port, regs_nxt_27_27_port, 
      regs_nxt_27_26_port, regs_nxt_27_25_port, regs_nxt_27_24_port, 
      regs_nxt_27_23_port, regs_nxt_27_22_port, regs_nxt_27_21_port, 
      regs_nxt_27_20_port, regs_nxt_27_19_port, regs_nxt_27_18_port, 
      regs_nxt_27_17_port, regs_nxt_27_16_port, regs_nxt_27_15_port, 
      regs_nxt_27_14_port, regs_nxt_27_13_port, regs_nxt_27_12_port, 
      regs_nxt_27_11_port, regs_nxt_27_10_port, regs_nxt_27_9_port, 
      regs_nxt_27_8_port, regs_nxt_27_7_port, regs_nxt_27_6_port, 
      regs_nxt_27_5_port, regs_nxt_27_4_port, regs_nxt_27_3_port, 
      regs_nxt_27_2_port, regs_nxt_27_1_port, regs_nxt_27_0_port, 
      regs_nxt_28_31_port, regs_nxt_28_30_port, regs_nxt_28_29_port, 
      regs_nxt_28_28_port, regs_nxt_28_27_port, regs_nxt_28_26_port, 
      regs_nxt_28_25_port, regs_nxt_28_24_port, regs_nxt_28_23_port, 
      regs_nxt_28_22_port, regs_nxt_28_21_port, regs_nxt_28_20_port, 
      regs_nxt_28_19_port, regs_nxt_28_18_port, regs_nxt_28_17_port, 
      regs_nxt_28_16_port, regs_nxt_28_15_port, regs_nxt_28_14_port, 
      regs_nxt_28_13_port, regs_nxt_28_12_port, regs_nxt_28_11_port, 
      regs_nxt_28_10_port, regs_nxt_28_9_port, regs_nxt_28_8_port, 
      regs_nxt_28_7_port, regs_nxt_28_6_port, regs_nxt_28_5_port, 
      regs_nxt_28_4_port, regs_nxt_28_3_port, regs_nxt_28_2_port, 
      regs_nxt_28_1_port, regs_nxt_28_0_port, regs_nxt_29_31_port, 
      regs_nxt_29_30_port, regs_nxt_29_29_port, regs_nxt_29_28_port, 
      regs_nxt_29_27_port, regs_nxt_29_26_port, regs_nxt_29_25_port, 
      regs_nxt_29_24_port, regs_nxt_29_23_port, regs_nxt_29_22_port, 
      regs_nxt_29_21_port, regs_nxt_29_20_port, regs_nxt_29_19_port, 
      regs_nxt_29_18_port, regs_nxt_29_17_port, regs_nxt_29_16_port, 
      regs_nxt_29_15_port, regs_nxt_29_14_port, regs_nxt_29_13_port, 
      regs_nxt_29_12_port, regs_nxt_29_11_port, regs_nxt_29_10_port, 
      regs_nxt_29_9_port, regs_nxt_29_8_port, regs_nxt_29_7_port, 
      regs_nxt_29_6_port, regs_nxt_29_5_port, regs_nxt_29_4_port, 
      regs_nxt_29_3_port, regs_nxt_29_2_port, regs_nxt_29_1_port, 
      regs_nxt_29_0_port, regs_nxt_30_31_port, regs_nxt_30_30_port, 
      regs_nxt_30_29_port, regs_nxt_30_28_port, regs_nxt_30_27_port, 
      regs_nxt_30_26_port, regs_nxt_30_25_port, regs_nxt_30_24_port, 
      regs_nxt_30_23_port, regs_nxt_30_22_port, regs_nxt_30_21_port, 
      regs_nxt_30_20_port, regs_nxt_30_19_port, regs_nxt_30_18_port, 
      regs_nxt_30_17_port, regs_nxt_30_16_port, regs_nxt_30_15_port, 
      regs_nxt_30_14_port, regs_nxt_30_13_port, regs_nxt_30_12_port, 
      regs_nxt_30_11_port, regs_nxt_30_10_port, regs_nxt_30_9_port, 
      regs_nxt_30_8_port, regs_nxt_30_7_port, regs_nxt_30_6_port, 
      regs_nxt_30_5_port, regs_nxt_30_4_port, regs_nxt_30_3_port, 
      regs_nxt_30_2_port, regs_nxt_30_1_port, regs_nxt_30_0_port, 
      regs_nxt_31_31_port, regs_nxt_31_30_port, regs_nxt_31_29_port, 
      regs_nxt_31_28_port, regs_nxt_31_27_port, regs_nxt_31_26_port, 
      regs_nxt_31_25_port, regs_nxt_31_24_port, regs_nxt_31_23_port, 
      regs_nxt_31_22_port, regs_nxt_31_21_port, regs_nxt_31_20_port, 
      regs_nxt_31_19_port, regs_nxt_31_18_port, regs_nxt_31_17_port, 
      regs_nxt_31_16_port, regs_nxt_31_15_port, regs_nxt_31_14_port, 
      regs_nxt_31_13_port, regs_nxt_31_12_port, regs_nxt_31_11_port, 
      regs_nxt_31_10_port, regs_nxt_31_9_port, regs_nxt_31_8_port, 
      regs_nxt_31_7_port, regs_nxt_31_6_port, regs_nxt_31_5_port, 
      regs_nxt_31_4_port, regs_nxt_31_3_port, regs_nxt_31_2_port, 
      regs_nxt_31_1_port, regs_nxt_31_0_port, N23, N24, N25, N26, N27, N28, N29
      , N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, 
      N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58
      , N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, 
      N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87
      , N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
      N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, 
      N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, 
      N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, 
      N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, 
      N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, 
      N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, 
      N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, 
      N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, 
      N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, 
      N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, 
      N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
      N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, 
      N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, 
      N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, 
      N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, 
      N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, 
      N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, 
      N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, 
      N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, 
      N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, 
      N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, 
      N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, 
      N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, 
      N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, 
      N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, 
      N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, 
      N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, 
      N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, 
      N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, 
      N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, 
      N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, 
      N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, 
      N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, 
      N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, 
      N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, 
      N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, 
      N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, 
      N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, 
      N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, 
      N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, 
      N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, 
      N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, 
      N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, 
      N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, 
      N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, 
      N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, 
      N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, 
      N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, 
      N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, 
      N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, 
      N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, 
      N714, N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, 
      N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, 
      N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, 
      N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, 
      N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, 
      N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, 
      N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, 
      N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, 
      N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, 
      N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, 
      N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, 
      N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, 
      N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, 
      N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, 
      N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, 
      N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, 
      N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, 
      N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, 
      N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, 
      N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, 
      N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, 
      N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, 
      N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, 
      N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
      N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, 
      N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, 
      N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, 
      N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, 
      N1042, N1043, N1044, N1045, N1046, N2166, N2199, N2231, N2263, N2295, 
      N2327, N2359, N2391, N2423, N2455, N2487, N2519, N2551, N2583, N2615, 
      N2647, N2679, N2711, N2743, N2775, N2807, N2839, N2871, N2903, N2935, 
      N2967, N2999, N3031, N3063, N3095, N3127, N3159, n2546, n2547, n2548, 
      n2550, n2551_port, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559
      , n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
      n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, 
      n2580, n2581, n2582, n2583_port, n2584, n2585, n2586, n2587, n2588, n2589
      , n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
      n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
      n2610, n2611, n2612, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
      n2645, n2646, n2647_port, n2648, n2649, n2650, n2651, n2652, n2653, n2654
      , n2655, n2656, n2657, n25179, n25180, n25181, n25182, n25183, n25184, 
      n25185, n25186, n25211, n25212, n25213, n25214, n25215, n25216, n25217, 
      n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, 
      n25227, n25228, n25229, n25230, n25236, n25237, n25238, n25239, n25240, 
      n25241, n25242, n25243, n25244, n25250, n25251, n25252, n25253, n25254, 
      n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, 
      n25264, n25265, n25266, n25267, n25268, n25269, n25291, n25292, n25293, 
      n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, 
      n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25434, 
      n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, 
      n25444, n25445, n25446, n25447, n25448, n25466, n25467, n25468, n25469, 
      n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, 
      n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25491, n25492, 
      n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, 
      n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, 
      n25511, n25512, n25513, n25514, n25515, n25516, n25532, n25533, n25534, 
      n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, 
      n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25557, 
      n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n635_port
      , n636_port, n637_port, n638_port, n639_port, n640_port, n641_port, 
      n642_port, n643_port, n644_port, n645_port, n646_port, n647_port, 
      n648_port, n649_port, n650_port, n651_port, n652_port, n653_port, 
      n654_port, n655_port, n656_port, n657_port, n658_port, n659_port, 
      n660_port, n661_port, n662_port, n663_port, n664_port, n665_port, 
      n666_port, n667_port, n668_port, n669_port, n670_port, n671_port, 
      n672_port, n673_port, n674_port, n675_port, n678_port, n679_port, 
      n680_port, n681_port, n682_port, n683_port, n684_port, n685_port, 
      n686_port, n687_port, n688_port, n689_port, n690_port, n691_port, 
      n692_port, n693_port, n694_port, n695_port, n696_port, n697_port, 
      n698_port, n699_port, n700_port, n701_port, n702_port, n703_port, 
      n704_port, n705_port, n706_port, n707_port, n708_port, n709_port, 
      n710_port, n711_port, n712_port, n713_port, n714_port, n715_port, 
      n716_port, n717_port, n718_port, n719_port, n720_port, n721_port, 
      n722_port, n723_port, n724_port, n725_port, n726_port, n727_port, 
      n728_port, n729_port, n730_port, n731_port, n732_port, n733_port, 
      n734_port, n735_port, n736_port, n737_port, n738_port, n739_port, 
      n740_port, n741_port, n742_port, n743_port, n744_port, n745_port, 
      n746_port, n747_port, n748_port, n749_port, n750_port, n751_port, 
      n752_port, n753_port, n754_port, n755_port, n756_port, n757_port, 
      n758_port, n759_port, n760_port, n761_port, n762_port, n763_port, 
      n764_port, n765_port, n766_port, n767_port, n768_port, n769_port, 
      n770_port, n771_port, n772_port, n773_port, n774_port, n775_port, 
      n776_port, n777_port, n778_port, n779_port, n780_port, n781_port, 
      n782_port, n783_port, n784_port, n785_port, n786_port, n787_port, 
      n788_port, n789_port, n790_port, n791_port, n792_port, n793_port, 
      n794_port, n795_port, n796_port, n797_port, n798_port, n799_port, 
      n800_port, n801_port, n802_port, n803_port, n804_port, n805_port, 
      n806_port, n807_port, n808_port, n809_port, n810_port, n811_port, 
      n812_port, n813_port, n814_port, n815_port, n816_port, n817_port, 
      n818_port, n819_port, n820_port, n821_port, n822_port, n823_port, 
      n824_port, n825_port, n826_port, n827_port, n828_port, n829_port, 
      n830_port, n831_port, n832_port, n833_port, n834_port, n835_port, 
      n836_port, n837_port, n838_port, n839_port, n840_port, n841_port, 
      n842_port, n843_port, n844_port, n845_port, n846_port, n847_port, 
      n848_port, n849_port, n850_port, n851_port, n852_port, n853_port, 
      n854_port, n855_port, n856_port, n857_port, n858_port, n859_port, 
      n860_port, n861_port, n862_port, n863_port, n864_port, n865_port, 
      n866_port, n867_port, n868_port, n869_port, n870_port, n871_port, 
      n872_port, n873_port, n874_port, n875_port, n876_port, n877_port, 
      n878_port, n879_port, n880_port, n881_port, n882_port, n883_port, 
      n884_port, n885_port, n886_port, n887_port, n888_port, n889_port, 
      n890_port, n891_port, n892_port, n893_port, n894_port, n895_port, 
      n896_port, n897_port, n898_port, n899_port, n900_port, n901_port, 
      n902_port, n903_port, n904_port, n905_port, n906_port, n907_port, 
      n908_port, n909_port, n910_port, n911_port, n912_port, n913_port, 
      n914_port, n915_port, n916_port, n917_port, n918_port, n919_port, 
      n920_port, n921_port, n922_port, n923_port, n924_port, n925_port, 
      n926_port, n927_port, n928_port, n929_port, n930_port, n931_port, 
      n932_port, n933_port, n934_port, n935_port, n936_port, n937_port, 
      n938_port, n939_port, n940_port, n941_port, n942_port, n943_port, 
      n944_port, n945_port, n946_port, n947_port, n948_port, n949_port, 
      n950_port, n951_port, n952_port, n953_port, n954_port, n955_port, 
      n956_port, n957_port, n958_port, n959_port, n960_port, n961_port, 
      n962_port, n963_port, n964_port, n965_port, n966_port, n967_port, 
      n968_port, n969_port, n970_port, n971_port, n972_port, n973_port, 
      n974_port, n975_port, n976_port, n977_port, n978_port, n979_port, 
      n980_port, n981_port, n982_port, n983_port, n984_port, n985_port, 
      n986_port, n987_port, n988_port, n989_port, n990_port, n991_port, 
      n992_port, n993_port, n994_port, n995_port, n996_port, n997_port, 
      n998_port, n999_port, n1000_port, n1001_port, n1002_port, n1003_port, 
      n1004_port, n1005_port, n1006_port, n1007_port, n1008_port, n1009_port, 
      n1010_port, n1011_port, n1012_port, n1013_port, n1014_port, n1015_port, 
      n1016_port, n1017_port, n1018_port, n1019_port, n1020_port, n1021_port, 
      n1022_port, n1023_port, n1024_port, n1025_port, n1026_port, n1027_port, 
      n1028_port, n1029_port, n1030_port, n1031_port, n1032_port, n1033_port, 
      n1034_port, n1035_port, n1036_port, n1037_port, n1038_port, n1039_port, 
      n1040_port, n1041_port, n1042_port, n1043_port, n1044_port, n1045_port, 
      n1046_port, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055
      , n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, 
      n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, 
      n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, 
      n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, 
      n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, 
      n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
      n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
      n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, 
      n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, 
      n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, 
      n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, 
      n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, 
      n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, 
      n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, 
      n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
      n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, 
      n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
      n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, 
      n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, 
      n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, 
      n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, 
      n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, 
      n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
      n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
      n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
      n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, 
      n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, 
      n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
      n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, 
      n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
      n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, 
      n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, 
      n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, 
      n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, 
      n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, 
      n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
      n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
      n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, 
      n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
      n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, 
      n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, 
      n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, 
      n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, 
      n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, 
      n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, 
      n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
      n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, 
      n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2079, 
      n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
      n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
      n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
      n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
      n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
      n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
      n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, 
      n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, 
      n2160, n2161, n2162, n2163, n2164, n2165, n2166_port, n2167, n2168, n2169
      , n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
      n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
      n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199_port
      , n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, 
      n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, 
      n2220, n2221, n2222, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295_port, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303
      , n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
      n2324, n2325, n2326, n2327_port, n2328, n2329, n2330, n2331, n2332, n2333
      , n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, 
      n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, 
      n2354, n2355, n2356, n2357, n2358, n2359_port, n2360, n2361, n2362, n2363
      , n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, 
      n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
      n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391_port, n2392, n2393
      , n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, 
      n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, 
      n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423_port
      , n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, 
      n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, 
      n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, 
      n2454, n2455_port, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463
      , n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, 
      n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, 
      n2484, n2485, n2486, n26327, n26328, n26329, n26330, n26331, n26332, 
      n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, 
      n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, 
      n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, 
      n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, 
      n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, 
      n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, 
      n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, 
      n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, 
      n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, 
      n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, 
      n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, 
      n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, 
      n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, 
      n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, 
      n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, 
      n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, 
      n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, 
      n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, 
      n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, 
      n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, 
      n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, 
      n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, 
      n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, 
      n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, 
      n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, 
      n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, 
      n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, 
      n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, 
      n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, 
      n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, 
      n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, 
      n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, 
      n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, 
      n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, 
      n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, 
      n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, 
      n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, 
      n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, 
      n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, 
      n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, 
      n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, 
      n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, 
      n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, 
      n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, 
      n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, 
      n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, 
      n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, 
      n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, 
      n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, 
      n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, 
      n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, 
      n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, 
      n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, 
      n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, 
      n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, 
      n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, 
      n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, 
      n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, 
      n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, 
      n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, 
      n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, 
      n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, 
      n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, 
      n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, 
      n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, 
      n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, 
      n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, 
      n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, 
      n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, 
      n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, 
      n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, 
      n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, 
      n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, 
      n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, 
      n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, 
      n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, 
      n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, 
      n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, 
      n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, 
      n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, 
      n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, 
      n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, 
      n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, 
      n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, 
      n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, 
      n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, 
      n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, 
      n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, 
      n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, 
      n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, 
      n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, 
      n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, 
      n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, 
      n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, 
      n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, 
      n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, 
      n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, 
      n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, 
      n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, 
      n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, 
      n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, 
      n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, 
      n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, 
      n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, 
      n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, 
      n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, 
      n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, 
      n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, 
      n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, 
      n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, 
      n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, 
      n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, 
      n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, 
      n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, 
      n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, 
      n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, 
      n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, 
      n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, 
      n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, 
      n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, 
      n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, 
      n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, 
      n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, 
      n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, 
      n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, 
      n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, 
      n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, 
      n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, 
      n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, 
      n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, 
      n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, 
      n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, 
      n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, 
      n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, 
      n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, 
      n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, 
      n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, 
      n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, 
      n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, 
      n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, 
      n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, 
      n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, 
      n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, 
      n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, 
      n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, 
      n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, 
      n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, 
      n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, 
      n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, 
      n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, 
      n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, 
      n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, 
      n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, 
      n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, 
      n27719, n27720, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626 : std_logic;

begin
   
   regs_nxt_reg_0_31_inst : DLH_X1 port map( G => n27469, D => n27373, Q => 
                           regs_nxt_0_31_port);
   regs_reg_0_31_inst : DFF_X1 port map( D => N1046, CK => clk, Q => n_1067, QN
                           => n26358);
   regs_nxt_reg_0_30_inst : DLH_X1 port map( G => n27469, D => n27379, Q => 
                           regs_nxt_0_30_port);
   regs_reg_0_30_inst : DFF_X1 port map( D => N1045, CK => clk, Q => n_1068, QN
                           => n26357);
   regs_nxt_reg_0_29_inst : DLH_X1 port map( G => n27468, D => n27385, Q => 
                           regs_nxt_0_29_port);
   regs_reg_0_29_inst : DFF_X1 port map( D => N1044, CK => clk, Q => n_1069, QN
                           => n26356);
   regs_nxt_reg_0_28_inst : DLH_X1 port map( G => n27468, D => n27391, Q => 
                           regs_nxt_0_28_port);
   regs_reg_0_28_inst : DFF_X1 port map( D => N1043, CK => clk, Q => n_1070, QN
                           => n26355);
   regs_nxt_reg_0_27_inst : DLH_X1 port map( G => n27471, D => n27397, Q => 
                           regs_nxt_0_27_port);
   regs_reg_0_27_inst : DFF_X1 port map( D => N1042, CK => clk, Q => n_1071, QN
                           => n26354);
   regs_nxt_reg_0_26_inst : DLH_X1 port map( G => n27470, D => n27403, Q => 
                           regs_nxt_0_26_port);
   regs_reg_0_26_inst : DFF_X1 port map( D => N1041, CK => clk, Q => n_1072, QN
                           => n26353);
   regs_nxt_reg_0_25_inst : DLH_X1 port map( G => n27471, D => n27409, Q => 
                           regs_nxt_0_25_port);
   regs_reg_0_25_inst : DFF_X1 port map( D => N1040, CK => clk, Q => n_1073, QN
                           => n26352);
   regs_nxt_reg_0_24_inst : DLH_X1 port map( G => n27470, D => n27415, Q => 
                           regs_nxt_0_24_port);
   regs_reg_0_24_inst : DFF_X1 port map( D => N1039, CK => clk, Q => n_1074, QN
                           => n26351);
   regs_nxt_reg_0_23_inst : DLH_X1 port map( G => n27470, D => n27421, Q => 
                           regs_nxt_0_23_port);
   regs_reg_0_23_inst : DFF_X1 port map( D => N1038, CK => clk, Q => n_1075, QN
                           => n26350);
   regs_nxt_reg_0_22_inst : DLH_X1 port map( G => n27470, D => n27427, Q => 
                           regs_nxt_0_22_port);
   regs_reg_0_22_inst : DFF_X1 port map( D => N1037, CK => clk, Q => n_1076, QN
                           => n26349);
   regs_nxt_reg_0_21_inst : DLH_X1 port map( G => n27468, D => n27433, Q => 
                           regs_nxt_0_21_port);
   regs_reg_0_21_inst : DFF_X1 port map( D => N1036, CK => clk, Q => n_1077, QN
                           => n26348);
   regs_nxt_reg_0_20_inst : DLH_X1 port map( G => n27468, D => n27283, Q => 
                           regs_nxt_0_20_port);
   regs_reg_0_20_inst : DFF_X1 port map( D => N1035, CK => clk, Q => n_1078, QN
                           => n26347);
   regs_nxt_reg_0_19_inst : DLH_X1 port map( G => n27468, D => n27289, Q => 
                           regs_nxt_0_19_port);
   regs_reg_0_19_inst : DFF_X1 port map( D => N1034, CK => clk, Q => n_1079, QN
                           => n26346);
   regs_nxt_reg_0_18_inst : DLH_X1 port map( G => n27470, D => n27295, Q => 
                           regs_nxt_0_18_port);
   regs_reg_0_18_inst : DFF_X1 port map( D => N1033, CK => clk, Q => n_1080, QN
                           => n26345);
   regs_nxt_reg_0_17_inst : DLH_X1 port map( G => n27468, D => n27301, Q => 
                           regs_nxt_0_17_port);
   regs_reg_0_17_inst : DFF_X1 port map( D => N1032, CK => clk, Q => n_1081, QN
                           => n26344);
   regs_nxt_reg_0_16_inst : DLH_X1 port map( G => n27470, D => n27307, Q => 
                           regs_nxt_0_16_port);
   regs_reg_0_16_inst : DFF_X1 port map( D => N1031, CK => clk, Q => n_1082, QN
                           => n26343);
   regs_nxt_reg_0_15_inst : DLH_X1 port map( G => n27468, D => n27313, Q => 
                           regs_nxt_0_15_port);
   regs_reg_0_15_inst : DFF_X1 port map( D => N1030, CK => clk, Q => n_1083, QN
                           => n26342);
   regs_nxt_reg_0_14_inst : DLH_X1 port map( G => n27470, D => n27319, Q => 
                           regs_nxt_0_14_port);
   regs_reg_0_14_inst : DFF_X1 port map( D => N1029, CK => clk, Q => n_1084, QN
                           => n26341);
   regs_nxt_reg_0_13_inst : DLH_X1 port map( G => n27470, D => n27325, Q => 
                           regs_nxt_0_13_port);
   regs_reg_0_13_inst : DFF_X1 port map( D => N1028, CK => clk, Q => n_1085, QN
                           => n26340);
   regs_nxt_reg_0_12_inst : DLH_X1 port map( G => n27470, D => n27331, Q => 
                           regs_nxt_0_12_port);
   regs_reg_0_12_inst : DFF_X1 port map( D => N1027, CK => clk, Q => n_1086, QN
                           => n26339);
   regs_nxt_reg_0_11_inst : DLH_X1 port map( G => n27468, D => n27337, Q => 
                           regs_nxt_0_11_port);
   regs_reg_0_11_inst : DFF_X1 port map( D => N1026, CK => clk, Q => n_1087, QN
                           => n26338);
   regs_nxt_reg_0_10_inst : DLH_X1 port map( G => n27468, D => n27343, Q => 
                           regs_nxt_0_10_port);
   regs_reg_0_10_inst : DFF_X1 port map( D => N1025, CK => clk, Q => n_1088, QN
                           => n26337);
   regs_nxt_reg_0_9_inst : DLH_X1 port map( G => n27469, D => n27349, Q => 
                           regs_nxt_0_9_port);
   regs_reg_0_9_inst : DFF_X1 port map( D => N1024, CK => clk, Q => n_1089, QN 
                           => n26336);
   regs_nxt_reg_0_8_inst : DLH_X1 port map( G => n27469, D => n27355, Q => 
                           regs_nxt_0_8_port);
   regs_reg_0_8_inst : DFF_X1 port map( D => N1023, CK => clk, Q => n_1090, QN 
                           => n26335);
   regs_nxt_reg_0_7_inst : DLH_X1 port map( G => n27469, D => n27361, Q => 
                           regs_nxt_0_7_port);
   regs_reg_0_7_inst : DFF_X1 port map( D => N1022, CK => clk, Q => n_1091, QN 
                           => n26334);
   regs_nxt_reg_0_6_inst : DLH_X1 port map( G => n27469, D => n27367, Q => 
                           regs_nxt_0_6_port);
   regs_reg_0_6_inst : DFF_X1 port map( D => N1021, CK => clk, Q => n_1092, QN 
                           => n26333);
   regs_nxt_reg_0_5_inst : DLH_X1 port map( G => n27469, D => n27277, Q => 
                           regs_nxt_0_5_port);
   regs_reg_0_5_inst : DFF_X1 port map( D => N1020, CK => clk, Q => n_1093, QN 
                           => n26332);
   regs_nxt_reg_0_4_inst : DLH_X1 port map( G => n27469, D => n27439, Q => 
                           regs_nxt_0_4_port);
   regs_reg_0_4_inst : DFF_X1 port map( D => N1019, CK => clk, Q => n_1094, QN 
                           => n26331);
   regs_nxt_reg_0_3_inst : DLH_X1 port map( G => n27470, D => n27445, Q => 
                           regs_nxt_0_3_port);
   regs_reg_0_3_inst : DFF_X1 port map( D => N1018, CK => clk, Q => n_1095, QN 
                           => n26330);
   regs_nxt_reg_0_2_inst : DLH_X1 port map( G => n27469, D => n27451, Q => 
                           regs_nxt_0_2_port);
   regs_reg_0_2_inst : DFF_X1 port map( D => N1017, CK => clk, Q => n_1096, QN 
                           => n26329);
   regs_nxt_reg_0_1_inst : DLH_X1 port map( G => n27468, D => n27457, Q => 
                           regs_nxt_0_1_port);
   regs_reg_0_1_inst : DFF_X1 port map( D => N1016, CK => clk, Q => n_1097, QN 
                           => n26328);
   regs_nxt_reg_0_0_inst : DLH_X1 port map( G => n27469, D => n27463, Q => 
                           regs_nxt_0_0_port);
   regs_reg_0_0_inst : DFF_X1 port map( D => N1015, CK => clk, Q => n_1098, QN 
                           => n26327);
   regs_nxt_reg_1_31_inst : DLH_X1 port map( G => n27476, D => n27373, Q => 
                           regs_nxt_1_31_port);
   regs_reg_1_31_inst : DFF_X1 port map( D => N1014, CK => clk, Q => n_1099, QN
                           => n26390);
   regs_nxt_reg_1_30_inst : DLH_X1 port map( G => n27476, D => n27379, Q => 
                           regs_nxt_1_30_port);
   regs_reg_1_30_inst : DFF_X1 port map( D => N1013, CK => clk, Q => n_1100, QN
                           => n26389);
   regs_nxt_reg_1_29_inst : DLH_X1 port map( G => n27475, D => n27385, Q => 
                           regs_nxt_1_29_port);
   regs_reg_1_29_inst : DFF_X1 port map( D => N1012, CK => clk, Q => n_1101, QN
                           => n26388);
   regs_nxt_reg_1_28_inst : DLH_X1 port map( G => n27475, D => n27391, Q => 
                           regs_nxt_1_28_port);
   regs_reg_1_28_inst : DFF_X1 port map( D => N1011, CK => clk, Q => n_1102, QN
                           => n26387);
   regs_nxt_reg_1_27_inst : DLH_X1 port map( G => n27478, D => n27397, Q => 
                           regs_nxt_1_27_port);
   regs_reg_1_27_inst : DFF_X1 port map( D => N1010, CK => clk, Q => n_1103, QN
                           => n26386);
   regs_nxt_reg_1_26_inst : DLH_X1 port map( G => n27477, D => n27403, Q => 
                           regs_nxt_1_26_port);
   regs_reg_1_26_inst : DFF_X1 port map( D => N1009, CK => clk, Q => n_1104, QN
                           => n26385);
   regs_nxt_reg_1_25_inst : DLH_X1 port map( G => n27478, D => n27409, Q => 
                           regs_nxt_1_25_port);
   regs_reg_1_25_inst : DFF_X1 port map( D => N1008, CK => clk, Q => n_1105, QN
                           => n26384);
   regs_nxt_reg_1_24_inst : DLH_X1 port map( G => n27477, D => n27415, Q => 
                           regs_nxt_1_24_port);
   regs_reg_1_24_inst : DFF_X1 port map( D => N1007, CK => clk, Q => n_1106, QN
                           => n26383);
   regs_nxt_reg_1_23_inst : DLH_X1 port map( G => n27477, D => n27421, Q => 
                           regs_nxt_1_23_port);
   regs_reg_1_23_inst : DFF_X1 port map( D => N1006, CK => clk, Q => n_1107, QN
                           => n26382);
   regs_nxt_reg_1_22_inst : DLH_X1 port map( G => n27477, D => n27427, Q => 
                           regs_nxt_1_22_port);
   regs_reg_1_22_inst : DFF_X1 port map( D => N1005, CK => clk, Q => n_1108, QN
                           => n26381);
   regs_nxt_reg_1_21_inst : DLH_X1 port map( G => n27475, D => n27433, Q => 
                           regs_nxt_1_21_port);
   regs_reg_1_21_inst : DFF_X1 port map( D => N1004, CK => clk, Q => n_1109, QN
                           => n26380);
   regs_nxt_reg_1_20_inst : DLH_X1 port map( G => n27475, D => n27283, Q => 
                           regs_nxt_1_20_port);
   regs_reg_1_20_inst : DFF_X1 port map( D => N1003, CK => clk, Q => n_1110, QN
                           => n26379);
   regs_nxt_reg_1_19_inst : DLH_X1 port map( G => n27475, D => n27289, Q => 
                           regs_nxt_1_19_port);
   regs_reg_1_19_inst : DFF_X1 port map( D => N1002, CK => clk, Q => n_1111, QN
                           => n26378);
   regs_nxt_reg_1_18_inst : DLH_X1 port map( G => n27477, D => n27295, Q => 
                           regs_nxt_1_18_port);
   regs_reg_1_18_inst : DFF_X1 port map( D => N1001, CK => clk, Q => n_1112, QN
                           => n26377);
   regs_nxt_reg_1_17_inst : DLH_X1 port map( G => n27475, D => n27301, Q => 
                           regs_nxt_1_17_port);
   regs_reg_1_17_inst : DFF_X1 port map( D => N1000, CK => clk, Q => n_1113, QN
                           => n26376);
   regs_nxt_reg_1_16_inst : DLH_X1 port map( G => n27477, D => n27307, Q => 
                           regs_nxt_1_16_port);
   regs_reg_1_16_inst : DFF_X1 port map( D => N999, CK => clk, Q => n_1114, QN 
                           => n26375);
   regs_nxt_reg_1_15_inst : DLH_X1 port map( G => n27475, D => n27313, Q => 
                           regs_nxt_1_15_port);
   regs_reg_1_15_inst : DFF_X1 port map( D => N998, CK => clk, Q => n_1115, QN 
                           => n26374);
   regs_nxt_reg_1_14_inst : DLH_X1 port map( G => n27477, D => n27319, Q => 
                           regs_nxt_1_14_port);
   regs_reg_1_14_inst : DFF_X1 port map( D => N997, CK => clk, Q => n_1116, QN 
                           => n26373);
   regs_nxt_reg_1_13_inst : DLH_X1 port map( G => n27477, D => n27325, Q => 
                           regs_nxt_1_13_port);
   regs_reg_1_13_inst : DFF_X1 port map( D => N996, CK => clk, Q => n_1117, QN 
                           => n26372);
   regs_nxt_reg_1_12_inst : DLH_X1 port map( G => n27477, D => n27331, Q => 
                           regs_nxt_1_12_port);
   regs_reg_1_12_inst : DFF_X1 port map( D => N995, CK => clk, Q => n_1118, QN 
                           => n26371);
   regs_nxt_reg_1_11_inst : DLH_X1 port map( G => n27475, D => n27337, Q => 
                           regs_nxt_1_11_port);
   regs_reg_1_11_inst : DFF_X1 port map( D => N994, CK => clk, Q => n_1119, QN 
                           => n26370);
   regs_nxt_reg_1_10_inst : DLH_X1 port map( G => n27475, D => n27343, Q => 
                           regs_nxt_1_10_port);
   regs_reg_1_10_inst : DFF_X1 port map( D => N993, CK => clk, Q => n_1120, QN 
                           => n26369);
   regs_nxt_reg_1_9_inst : DLH_X1 port map( G => n27476, D => n27349, Q => 
                           regs_nxt_1_9_port);
   regs_reg_1_9_inst : DFF_X1 port map( D => N992, CK => clk, Q => n_1121, QN 
                           => n26368);
   regs_nxt_reg_1_8_inst : DLH_X1 port map( G => n27476, D => n27355, Q => 
                           regs_nxt_1_8_port);
   regs_reg_1_8_inst : DFF_X1 port map( D => N991, CK => clk, Q => n_1122, QN 
                           => n26367);
   regs_nxt_reg_1_7_inst : DLH_X1 port map( G => n27476, D => n27361, Q => 
                           regs_nxt_1_7_port);
   regs_reg_1_7_inst : DFF_X1 port map( D => N990, CK => clk, Q => n_1123, QN 
                           => n26366);
   regs_nxt_reg_1_6_inst : DLH_X1 port map( G => n27476, D => n27367, Q => 
                           regs_nxt_1_6_port);
   regs_reg_1_6_inst : DFF_X1 port map( D => N989, CK => clk, Q => n_1124, QN 
                           => n26365);
   regs_nxt_reg_1_5_inst : DLH_X1 port map( G => n27476, D => n27277, Q => 
                           regs_nxt_1_5_port);
   regs_reg_1_5_inst : DFF_X1 port map( D => N988, CK => clk, Q => n_1125, QN 
                           => n26364);
   regs_nxt_reg_1_4_inst : DLH_X1 port map( G => n27476, D => n27439, Q => 
                           regs_nxt_1_4_port);
   regs_reg_1_4_inst : DFF_X1 port map( D => N987, CK => clk, Q => n_1126, QN 
                           => n26363);
   regs_nxt_reg_1_3_inst : DLH_X1 port map( G => n27477, D => n27445, Q => 
                           regs_nxt_1_3_port);
   regs_reg_1_3_inst : DFF_X1 port map( D => N986, CK => clk, Q => n_1127, QN 
                           => n26362);
   regs_nxt_reg_1_2_inst : DLH_X1 port map( G => n27476, D => n27451, Q => 
                           regs_nxt_1_2_port);
   regs_reg_1_2_inst : DFF_X1 port map( D => N985, CK => clk, Q => n_1128, QN 
                           => n26361);
   regs_nxt_reg_1_1_inst : DLH_X1 port map( G => n27475, D => n27457, Q => 
                           regs_nxt_1_1_port);
   regs_reg_1_1_inst : DFF_X1 port map( D => N984, CK => clk, Q => n_1129, QN 
                           => n26360);
   regs_nxt_reg_1_0_inst : DLH_X1 port map( G => n27476, D => n27463, Q => 
                           regs_nxt_1_0_port);
   regs_reg_1_0_inst : DFF_X1 port map( D => N983, CK => clk, Q => n_1130, QN 
                           => n26359);
   regs_nxt_reg_2_31_inst : DLH_X1 port map( G => n27483, D => n27372, Q => 
                           regs_nxt_2_31_port);
   regs_reg_2_31_inst : DFF_X1 port map( D => N982, CK => clk, Q => n2216, QN 
                           => n26572);
   regs_nxt_reg_2_30_inst : DLH_X1 port map( G => n27483, D => n27378, Q => 
                           regs_nxt_2_30_port);
   regs_reg_2_30_inst : DFF_X1 port map( D => N981, CK => clk, Q => n2209, QN 
                           => n26570);
   regs_nxt_reg_2_29_inst : DLH_X1 port map( G => n27482, D => n27384, Q => 
                           regs_nxt_2_29_port);
   regs_reg_2_29_inst : DFF_X1 port map( D => N980, CK => clk, Q => n2202, QN 
                           => n26568);
   regs_nxt_reg_2_28_inst : DLH_X1 port map( G => n27482, D => n27390, Q => 
                           regs_nxt_2_28_port);
   regs_reg_2_28_inst : DFF_X1 port map( D => N979, CK => clk, Q => n2195, QN 
                           => n26566);
   regs_nxt_reg_2_27_inst : DLH_X1 port map( G => n27485, D => n27396, Q => 
                           regs_nxt_2_27_port);
   regs_reg_2_27_inst : DFF_X1 port map( D => N978, CK => clk, Q => n2188, QN 
                           => n26564);
   regs_nxt_reg_2_26_inst : DLH_X1 port map( G => n27484, D => n27402, Q => 
                           regs_nxt_2_26_port);
   regs_reg_2_26_inst : DFF_X1 port map( D => N977, CK => clk, Q => n2181, QN 
                           => n26562);
   regs_nxt_reg_2_25_inst : DLH_X1 port map( G => n27485, D => n27408, Q => 
                           regs_nxt_2_25_port);
   regs_reg_2_25_inst : DFF_X1 port map( D => N976, CK => clk, Q => n2174, QN 
                           => n26560);
   regs_nxt_reg_2_24_inst : DLH_X1 port map( G => n27484, D => n27414, Q => 
                           regs_nxt_2_24_port);
   regs_reg_2_24_inst : DFF_X1 port map( D => N975, CK => clk, Q => n2167, QN 
                           => n26558);
   regs_nxt_reg_2_23_inst : DLH_X1 port map( G => n27484, D => n27420, Q => 
                           regs_nxt_2_23_port);
   regs_reg_2_23_inst : DFF_X1 port map( D => N974, CK => clk, Q => n2160, QN 
                           => n26556);
   regs_nxt_reg_2_22_inst : DLH_X1 port map( G => n27484, D => n27426, Q => 
                           regs_nxt_2_22_port);
   regs_reg_2_22_inst : DFF_X1 port map( D => N973, CK => clk, Q => n2153, QN 
                           => n26554);
   regs_nxt_reg_2_21_inst : DLH_X1 port map( G => n27482, D => n27432, Q => 
                           regs_nxt_2_21_port);
   regs_reg_2_21_inst : DFF_X1 port map( D => N972, CK => clk, Q => n2146, QN 
                           => n26552);
   regs_nxt_reg_2_20_inst : DLH_X1 port map( G => n27482, D => n27282, Q => 
                           regs_nxt_2_20_port);
   regs_reg_2_20_inst : DFF_X1 port map( D => N971, CK => clk, Q => n2139, QN 
                           => n26550);
   regs_nxt_reg_2_19_inst : DLH_X1 port map( G => n27482, D => n27288, Q => 
                           regs_nxt_2_19_port);
   regs_reg_2_19_inst : DFF_X1 port map( D => N970, CK => clk, Q => n_1131, QN 
                           => n25551);
   regs_nxt_reg_2_18_inst : DLH_X1 port map( G => n27484, D => n27294, Q => 
                           regs_nxt_2_18_port);
   regs_reg_2_18_inst : DFF_X1 port map( D => N969, CK => clk, Q => n_1132, QN 
                           => n25550);
   regs_nxt_reg_2_17_inst : DLH_X1 port map( G => n27482, D => n27300, Q => 
                           regs_nxt_2_17_port);
   regs_reg_2_17_inst : DFF_X1 port map( D => N968, CK => clk, Q => n_1133, QN 
                           => n25549);
   regs_nxt_reg_2_16_inst : DLH_X1 port map( G => n27484, D => n27306, Q => 
                           regs_nxt_2_16_port);
   regs_reg_2_16_inst : DFF_X1 port map( D => N967, CK => clk, Q => n_1134, QN 
                           => n25548);
   regs_nxt_reg_2_15_inst : DLH_X1 port map( G => n27482, D => n27312, Q => 
                           regs_nxt_2_15_port);
   regs_reg_2_15_inst : DFF_X1 port map( D => N966, CK => clk, Q => n_1135, QN 
                           => n25547);
   regs_nxt_reg_2_14_inst : DLH_X1 port map( G => n27484, D => n27318, Q => 
                           regs_nxt_2_14_port);
   regs_reg_2_14_inst : DFF_X1 port map( D => N965, CK => clk, Q => n_1136, QN 
                           => n25546);
   regs_nxt_reg_2_13_inst : DLH_X1 port map( G => n27484, D => n27324, Q => 
                           regs_nxt_2_13_port);
   regs_reg_2_13_inst : DFF_X1 port map( D => N964, CK => clk, Q => n_1137, QN 
                           => n25545);
   regs_nxt_reg_2_12_inst : DLH_X1 port map( G => n27484, D => n27330, Q => 
                           regs_nxt_2_12_port);
   regs_reg_2_12_inst : DFF_X1 port map( D => N963, CK => clk, Q => n_1138, QN 
                           => n25544);
   regs_nxt_reg_2_11_inst : DLH_X1 port map( G => n27482, D => n27336, Q => 
                           regs_nxt_2_11_port);
   regs_reg_2_11_inst : DFF_X1 port map( D => N962, CK => clk, Q => n_1139, QN 
                           => n25543);
   regs_nxt_reg_2_10_inst : DLH_X1 port map( G => n27482, D => n27342, Q => 
                           regs_nxt_2_10_port);
   regs_reg_2_10_inst : DFF_X1 port map( D => N961, CK => clk, Q => n_1140, QN 
                           => n25542);
   regs_nxt_reg_2_9_inst : DLH_X1 port map( G => n27483, D => n27348, Q => 
                           regs_nxt_2_9_port);
   regs_reg_2_9_inst : DFF_X1 port map( D => N960, CK => clk, Q => n_1141, QN 
                           => n25541);
   regs_nxt_reg_2_8_inst : DLH_X1 port map( G => n27483, D => n27354, Q => 
                           regs_nxt_2_8_port);
   regs_reg_2_8_inst : DFF_X1 port map( D => N959, CK => clk, Q => n_1142, QN 
                           => n25540);
   regs_nxt_reg_2_7_inst : DLH_X1 port map( G => n27483, D => n27360, Q => 
                           regs_nxt_2_7_port);
   regs_reg_2_7_inst : DFF_X1 port map( D => N958, CK => clk, Q => n_1143, QN 
                           => n25539);
   regs_nxt_reg_2_6_inst : DLH_X1 port map( G => n27483, D => n27366, Q => 
                           regs_nxt_2_6_port);
   regs_reg_2_6_inst : DFF_X1 port map( D => N957, CK => clk, Q => n_1144, QN 
                           => n25538);
   regs_nxt_reg_2_5_inst : DLH_X1 port map( G => n27483, D => n27276, Q => 
                           regs_nxt_2_5_port);
   regs_reg_2_5_inst : DFF_X1 port map( D => N956, CK => clk, Q => n_1145, QN 
                           => n25537);
   regs_nxt_reg_2_4_inst : DLH_X1 port map( G => n27483, D => n27438, Q => 
                           regs_nxt_2_4_port);
   regs_reg_2_4_inst : DFF_X1 port map( D => N955, CK => clk, Q => n_1146, QN 
                           => n25536);
   regs_nxt_reg_2_3_inst : DLH_X1 port map( G => n27484, D => n27444, Q => 
                           regs_nxt_2_3_port);
   regs_reg_2_3_inst : DFF_X1 port map( D => N954, CK => clk, Q => n_1147, QN 
                           => n25535);
   regs_nxt_reg_2_2_inst : DLH_X1 port map( G => n27483, D => n27450, Q => 
                           regs_nxt_2_2_port);
   regs_reg_2_2_inst : DFF_X1 port map( D => N953, CK => clk, Q => n_1148, QN 
                           => n25534);
   regs_nxt_reg_2_1_inst : DLH_X1 port map( G => n27482, D => n27456, Q => 
                           regs_nxt_2_1_port);
   regs_reg_2_1_inst : DFF_X1 port map( D => N952, CK => clk, Q => n_1149, QN 
                           => n25533);
   regs_nxt_reg_2_0_inst : DLH_X1 port map( G => n27483, D => n27462, Q => 
                           regs_nxt_2_0_port);
   regs_reg_2_0_inst : DFF_X1 port map( D => N951, CK => clk, Q => n_1150, QN 
                           => n25532);
   regs_nxt_reg_3_31_inst : DLH_X1 port map( G => n27490, D => n27374, Q => 
                           regs_nxt_3_31_port);
   regs_reg_3_31_inst : DFF_X1 port map( D => N950, CK => clk, Q => n25499, QN 
                           => n_1151);
   regs_nxt_reg_3_30_inst : DLH_X1 port map( G => n27490, D => n27380, Q => 
                           regs_nxt_3_30_port);
   regs_reg_3_30_inst : DFF_X1 port map( D => N949, CK => clk, Q => n25498, QN 
                           => n_1152);
   regs_nxt_reg_3_29_inst : DLH_X1 port map( G => n27489, D => n27386, Q => 
                           regs_nxt_3_29_port);
   regs_reg_3_29_inst : DFF_X1 port map( D => N948, CK => clk, Q => n25497, QN 
                           => n_1153);
   regs_nxt_reg_3_28_inst : DLH_X1 port map( G => n27489, D => n27392, Q => 
                           regs_nxt_3_28_port);
   regs_reg_3_28_inst : DFF_X1 port map( D => N947, CK => clk, Q => n25496, QN 
                           => n_1154);
   regs_nxt_reg_3_27_inst : DLH_X1 port map( G => n27492, D => n27398, Q => 
                           regs_nxt_3_27_port);
   regs_reg_3_27_inst : DFF_X1 port map( D => N946, CK => clk, Q => n25495, QN 
                           => n_1155);
   regs_nxt_reg_3_26_inst : DLH_X1 port map( G => n27491, D => n27404, Q => 
                           regs_nxt_3_26_port);
   regs_reg_3_26_inst : DFF_X1 port map( D => N945, CK => clk, Q => n25494, QN 
                           => n_1156);
   regs_nxt_reg_3_25_inst : DLH_X1 port map( G => n27492, D => n27410, Q => 
                           regs_nxt_3_25_port);
   regs_reg_3_25_inst : DFF_X1 port map( D => N944, CK => clk, Q => n25493, QN 
                           => n_1157);
   regs_nxt_reg_3_24_inst : DLH_X1 port map( G => n27491, D => n27416, Q => 
                           regs_nxt_3_24_port);
   regs_reg_3_24_inst : DFF_X1 port map( D => N943, CK => clk, Q => n25492, QN 
                           => n_1158);
   regs_nxt_reg_3_23_inst : DLH_X1 port map( G => n27491, D => n27422, Q => 
                           regs_nxt_3_23_port);
   regs_reg_3_23_inst : DFF_X1 port map( D => N942, CK => clk, Q => n25491, QN 
                           => n_1159);
   regs_nxt_reg_3_22_inst : DLH_X1 port map( G => n27491, D => n27428, Q => 
                           regs_nxt_3_22_port);
   regs_reg_3_22_inst : DFF_X1 port map( D => N941, CK => clk, Q => n26413, QN 
                           => n2357);
   regs_nxt_reg_3_21_inst : DLH_X1 port map( G => n27489, D => n27434, Q => 
                           regs_nxt_3_21_port);
   regs_reg_3_21_inst : DFF_X1 port map( D => N940, CK => clk, Q => n26412, QN 
                           => n2353);
   regs_nxt_reg_3_20_inst : DLH_X1 port map( G => n27489, D => n27284, Q => 
                           regs_nxt_3_20_port);
   regs_reg_3_20_inst : DFF_X1 port map( D => N939, CK => clk, Q => n26411, QN 
                           => n2349);
   regs_nxt_reg_3_19_inst : DLH_X1 port map( G => n27489, D => n27290, Q => 
                           regs_nxt_3_19_port);
   regs_reg_3_19_inst : DFF_X1 port map( D => N938, CK => clk, Q => n26410, QN 
                           => n2345);
   regs_nxt_reg_3_18_inst : DLH_X1 port map( G => n27491, D => n27296, Q => 
                           regs_nxt_3_18_port);
   regs_reg_3_18_inst : DFF_X1 port map( D => N937, CK => clk, Q => n26409, QN 
                           => n2341);
   regs_nxt_reg_3_17_inst : DLH_X1 port map( G => n27489, D => n27302, Q => 
                           regs_nxt_3_17_port);
   regs_reg_3_17_inst : DFF_X1 port map( D => N936, CK => clk, Q => n26408, QN 
                           => n2337);
   regs_nxt_reg_3_16_inst : DLH_X1 port map( G => n27491, D => n27308, Q => 
                           regs_nxt_3_16_port);
   regs_reg_3_16_inst : DFF_X1 port map( D => N935, CK => clk, Q => n26407, QN 
                           => n2333);
   regs_nxt_reg_3_15_inst : DLH_X1 port map( G => n27489, D => n27314, Q => 
                           regs_nxt_3_15_port);
   regs_reg_3_15_inst : DFF_X1 port map( D => N934, CK => clk, Q => n26406, QN 
                           => n2329);
   regs_nxt_reg_3_14_inst : DLH_X1 port map( G => n27491, D => n27320, Q => 
                           regs_nxt_3_14_port);
   regs_reg_3_14_inst : DFF_X1 port map( D => N933, CK => clk, Q => n26405, QN 
                           => n2325);
   regs_nxt_reg_3_13_inst : DLH_X1 port map( G => n27491, D => n27326, Q => 
                           regs_nxt_3_13_port);
   regs_reg_3_13_inst : DFF_X1 port map( D => N932, CK => clk, Q => n26404, QN 
                           => n2321);
   regs_nxt_reg_3_12_inst : DLH_X1 port map( G => n27491, D => n27332, Q => 
                           regs_nxt_3_12_port);
   regs_reg_3_12_inst : DFF_X1 port map( D => N931, CK => clk, Q => n26403, QN 
                           => n2317);
   regs_nxt_reg_3_11_inst : DLH_X1 port map( G => n27489, D => n27338, Q => 
                           regs_nxt_3_11_port);
   regs_reg_3_11_inst : DFF_X1 port map( D => N930, CK => clk, Q => n26402, QN 
                           => n2313);
   regs_nxt_reg_3_10_inst : DLH_X1 port map( G => n27489, D => n27344, Q => 
                           regs_nxt_3_10_port);
   regs_reg_3_10_inst : DFF_X1 port map( D => N929, CK => clk, Q => n26401, QN 
                           => n2309);
   regs_nxt_reg_3_9_inst : DLH_X1 port map( G => n27490, D => n27350, Q => 
                           regs_nxt_3_9_port);
   regs_reg_3_9_inst : DFF_X1 port map( D => N928, CK => clk, Q => n26400, QN 
                           => n2305);
   regs_nxt_reg_3_8_inst : DLH_X1 port map( G => n27490, D => n27356, Q => 
                           regs_nxt_3_8_port);
   regs_reg_3_8_inst : DFF_X1 port map( D => N927, CK => clk, Q => n26399, QN 
                           => n2301);
   regs_nxt_reg_3_7_inst : DLH_X1 port map( G => n27490, D => n27362, Q => 
                           regs_nxt_3_7_port);
   regs_reg_3_7_inst : DFF_X1 port map( D => N926, CK => clk, Q => n26398, QN 
                           => n2297);
   regs_nxt_reg_3_6_inst : DLH_X1 port map( G => n27490, D => n27368, Q => 
                           regs_nxt_3_6_port);
   regs_reg_3_6_inst : DFF_X1 port map( D => N925, CK => clk, Q => n26397, QN 
                           => n2293);
   regs_nxt_reg_3_5_inst : DLH_X1 port map( G => n27490, D => n27278, Q => 
                           regs_nxt_3_5_port);
   regs_reg_3_5_inst : DFF_X1 port map( D => N924, CK => clk, Q => n26396, QN 
                           => n2289);
   regs_nxt_reg_3_4_inst : DLH_X1 port map( G => n27490, D => n27440, Q => 
                           regs_nxt_3_4_port);
   regs_reg_3_4_inst : DFF_X1 port map( D => N923, CK => clk, Q => n26395, QN 
                           => n2657);
   regs_nxt_reg_3_3_inst : DLH_X1 port map( G => n27491, D => n27446, Q => 
                           regs_nxt_3_3_port);
   regs_reg_3_3_inst : DFF_X1 port map( D => N922, CK => clk, Q => n26394, QN 
                           => n2655);
   regs_nxt_reg_3_2_inst : DLH_X1 port map( G => n27490, D => n27452, Q => 
                           regs_nxt_3_2_port);
   regs_reg_3_2_inst : DFF_X1 port map( D => N921, CK => clk, Q => n26393, QN 
                           => n2653);
   regs_nxt_reg_3_1_inst : DLH_X1 port map( G => n27489, D => n27458, Q => 
                           regs_nxt_3_1_port);
   regs_reg_3_1_inst : DFF_X1 port map( D => N920, CK => clk, Q => n26392, QN 
                           => n2651);
   regs_nxt_reg_3_0_inst : DLH_X1 port map( G => n27490, D => n27464, Q => 
                           regs_nxt_3_0_port);
   regs_reg_3_0_inst : DFF_X1 port map( D => N919, CK => clk, Q => n26391, QN 
                           => n2649);
   regs_nxt_reg_4_31_inst : DLH_X1 port map( G => n27497, D => n27372, Q => 
                           regs_nxt_4_31_port);
   regs_reg_4_31_inst : DFF_X1 port map( D => N918, CK => clk, Q => n_1160, QN 
                           => n25565);
   regs_nxt_reg_4_30_inst : DLH_X1 port map( G => n27497, D => n27378, Q => 
                           regs_nxt_4_30_port);
   regs_reg_4_30_inst : DFF_X1 port map( D => N917, CK => clk, Q => n_1161, QN 
                           => n25564);
   regs_nxt_reg_4_29_inst : DLH_X1 port map( G => n27496, D => n27384, Q => 
                           regs_nxt_4_29_port);
   regs_reg_4_29_inst : DFF_X1 port map( D => N916, CK => clk, Q => n_1162, QN 
                           => n25563);
   regs_nxt_reg_4_28_inst : DLH_X1 port map( G => n27496, D => n27390, Q => 
                           regs_nxt_4_28_port);
   regs_reg_4_28_inst : DFF_X1 port map( D => N915, CK => clk, Q => n_1163, QN 
                           => n25562);
   regs_nxt_reg_4_27_inst : DLH_X1 port map( G => n27499, D => n27396, Q => 
                           regs_nxt_4_27_port);
   regs_reg_4_27_inst : DFF_X1 port map( D => N914, CK => clk, Q => n_1164, QN 
                           => n25561);
   regs_nxt_reg_4_26_inst : DLH_X1 port map( G => n27498, D => n27402, Q => 
                           regs_nxt_4_26_port);
   regs_reg_4_26_inst : DFF_X1 port map( D => N913, CK => clk, Q => n_1165, QN 
                           => n25560);
   regs_nxt_reg_4_25_inst : DLH_X1 port map( G => n27499, D => n27408, Q => 
                           regs_nxt_4_25_port);
   regs_reg_4_25_inst : DFF_X1 port map( D => N912, CK => clk, Q => n_1166, QN 
                           => n25559);
   regs_nxt_reg_4_24_inst : DLH_X1 port map( G => n27498, D => n27414, Q => 
                           regs_nxt_4_24_port);
   regs_reg_4_24_inst : DFF_X1 port map( D => N911, CK => clk, Q => n_1167, QN 
                           => n25558);
   regs_nxt_reg_4_23_inst : DLH_X1 port map( G => n27498, D => n27420, Q => 
                           regs_nxt_4_23_port);
   regs_reg_4_23_inst : DFF_X1 port map( D => N910, CK => clk, Q => n_1168, QN 
                           => n25557);
   regs_nxt_reg_4_22_inst : DLH_X1 port map( G => n27498, D => n27426, Q => 
                           regs_nxt_4_22_port);
   regs_reg_4_22_inst : DFF_X1 port map( D => N909, CK => clk, Q => n2355, QN 
                           => n26497);
   regs_nxt_reg_4_21_inst : DLH_X1 port map( G => n27496, D => n27432, Q => 
                           regs_nxt_4_21_port);
   regs_reg_4_21_inst : DFF_X1 port map( D => N908, CK => clk, Q => n2351, QN 
                           => n26496);
   regs_nxt_reg_4_20_inst : DLH_X1 port map( G => n27496, D => n27282, Q => 
                           regs_nxt_4_20_port);
   regs_reg_4_20_inst : DFF_X1 port map( D => N907, CK => clk, Q => n2347, QN 
                           => n26495);
   regs_nxt_reg_4_19_inst : DLH_X1 port map( G => n27496, D => n27288, Q => 
                           regs_nxt_4_19_port);
   regs_reg_4_19_inst : DFF_X1 port map( D => N906, CK => clk, Q => n2343, QN 
                           => n26494);
   regs_nxt_reg_4_18_inst : DLH_X1 port map( G => n27498, D => n27294, Q => 
                           regs_nxt_4_18_port);
   regs_reg_4_18_inst : DFF_X1 port map( D => N905, CK => clk, Q => n2339, QN 
                           => n26493);
   regs_nxt_reg_4_17_inst : DLH_X1 port map( G => n27496, D => n27300, Q => 
                           regs_nxt_4_17_port);
   regs_reg_4_17_inst : DFF_X1 port map( D => N904, CK => clk, Q => n2335, QN 
                           => n26492);
   regs_nxt_reg_4_16_inst : DLH_X1 port map( G => n27498, D => n27306, Q => 
                           regs_nxt_4_16_port);
   regs_reg_4_16_inst : DFF_X1 port map( D => N903, CK => clk, Q => n2331, QN 
                           => n26491);
   regs_nxt_reg_4_15_inst : DLH_X1 port map( G => n27496, D => n27312, Q => 
                           regs_nxt_4_15_port);
   regs_reg_4_15_inst : DFF_X1 port map( D => N902, CK => clk, Q => n2327_port,
                           QN => n26490);
   regs_nxt_reg_4_14_inst : DLH_X1 port map( G => n27498, D => n27318, Q => 
                           regs_nxt_4_14_port);
   regs_reg_4_14_inst : DFF_X1 port map( D => N901, CK => clk, Q => n2323, QN 
                           => n26489);
   regs_nxt_reg_4_13_inst : DLH_X1 port map( G => n27498, D => n27324, Q => 
                           regs_nxt_4_13_port);
   regs_reg_4_13_inst : DFF_X1 port map( D => N900, CK => clk, Q => n2319, QN 
                           => n26488);
   regs_nxt_reg_4_12_inst : DLH_X1 port map( G => n27498, D => n27330, Q => 
                           regs_nxt_4_12_port);
   regs_reg_4_12_inst : DFF_X1 port map( D => N899, CK => clk, Q => n2315, QN 
                           => n26487);
   regs_nxt_reg_4_11_inst : DLH_X1 port map( G => n27496, D => n27336, Q => 
                           regs_nxt_4_11_port);
   regs_reg_4_11_inst : DFF_X1 port map( D => N898, CK => clk, Q => n2311, QN 
                           => n26486);
   regs_nxt_reg_4_10_inst : DLH_X1 port map( G => n27496, D => n27342, Q => 
                           regs_nxt_4_10_port);
   regs_reg_4_10_inst : DFF_X1 port map( D => N897, CK => clk, Q => n2307, QN 
                           => n26485);
   regs_nxt_reg_4_9_inst : DLH_X1 port map( G => n27497, D => n27348, Q => 
                           regs_nxt_4_9_port);
   regs_reg_4_9_inst : DFF_X1 port map( D => N896, CK => clk, Q => n2303, QN =>
                           n26484);
   regs_nxt_reg_4_8_inst : DLH_X1 port map( G => n27497, D => n27354, Q => 
                           regs_nxt_4_8_port);
   regs_reg_4_8_inst : DFF_X1 port map( D => N895, CK => clk, Q => n2299, QN =>
                           n26483);
   regs_nxt_reg_4_7_inst : DLH_X1 port map( G => n27497, D => n27360, Q => 
                           regs_nxt_4_7_port);
   regs_reg_4_7_inst : DFF_X1 port map( D => N894, CK => clk, Q => n2295_port, 
                           QN => n26482);
   regs_nxt_reg_4_6_inst : DLH_X1 port map( G => n27497, D => n27366, Q => 
                           regs_nxt_4_6_port);
   regs_reg_4_6_inst : DFF_X1 port map( D => N893, CK => clk, Q => n2291, QN =>
                           n26481);
   regs_nxt_reg_4_5_inst : DLH_X1 port map( G => n27497, D => n27276, Q => 
                           regs_nxt_4_5_port);
   regs_reg_4_5_inst : DFF_X1 port map( D => N892, CK => clk, Q => n2287, QN =>
                           n26480);
   regs_nxt_reg_4_4_inst : DLH_X1 port map( G => n27497, D => n27438, Q => 
                           regs_nxt_4_4_port);
   regs_reg_4_4_inst : DFF_X1 port map( D => N891, CK => clk, Q => n2646, QN =>
                           n26479);
   regs_nxt_reg_4_3_inst : DLH_X1 port map( G => n27498, D => n27444, Q => 
                           regs_nxt_4_3_port);
   regs_reg_4_3_inst : DFF_X1 port map( D => N890, CK => clk, Q => n2644, QN =>
                           n26478);
   regs_nxt_reg_4_2_inst : DLH_X1 port map( G => n27497, D => n27450, Q => 
                           regs_nxt_4_2_port);
   regs_reg_4_2_inst : DFF_X1 port map( D => N889, CK => clk, Q => n2642, QN =>
                           n26477);
   regs_nxt_reg_4_1_inst : DLH_X1 port map( G => n27496, D => n27456, Q => 
                           regs_nxt_4_1_port);
   regs_reg_4_1_inst : DFF_X1 port map( D => N888, CK => clk, Q => n2640, QN =>
                           n26476);
   regs_nxt_reg_4_0_inst : DLH_X1 port map( G => n27497, D => n27462, Q => 
                           regs_nxt_4_0_port);
   regs_reg_4_0_inst : DFF_X1 port map( D => N887, CK => clk, Q => n2638, QN =>
                           n26475);
   regs_nxt_reg_5_31_inst : DLH_X1 port map( G => n27504, D => n27375, Q => 
                           regs_nxt_5_31_port);
   regs_reg_5_31_inst : DFF_X1 port map( D => N886, CK => clk, Q => 
                           regs_5_31_port, QN => n_1169);
   regs_nxt_reg_5_30_inst : DLH_X1 port map( G => n27504, D => n27381, Q => 
                           regs_nxt_5_30_port);
   regs_reg_5_30_inst : DFF_X1 port map( D => N885, CK => clk, Q => 
                           regs_5_30_port, QN => n_1170);
   regs_nxt_reg_5_29_inst : DLH_X1 port map( G => n27503, D => n27387, Q => 
                           regs_nxt_5_29_port);
   regs_reg_5_29_inst : DFF_X1 port map( D => N884, CK => clk, Q => 
                           regs_5_29_port, QN => n_1171);
   regs_nxt_reg_5_28_inst : DLH_X1 port map( G => n27503, D => n27393, Q => 
                           regs_nxt_5_28_port);
   regs_reg_5_28_inst : DFF_X1 port map( D => N883, CK => clk, Q => 
                           regs_5_28_port, QN => n_1172);
   regs_nxt_reg_5_27_inst : DLH_X1 port map( G => n27506, D => n27399, Q => 
                           regs_nxt_5_27_port);
   regs_reg_5_27_inst : DFF_X1 port map( D => N882, CK => clk, Q => 
                           regs_5_27_port, QN => n_1173);
   regs_nxt_reg_5_26_inst : DLH_X1 port map( G => n27505, D => n27405, Q => 
                           regs_nxt_5_26_port);
   regs_reg_5_26_inst : DFF_X1 port map( D => N881, CK => clk, Q => 
                           regs_5_26_port, QN => n_1174);
   regs_nxt_reg_5_25_inst : DLH_X1 port map( G => n27506, D => n27411, Q => 
                           regs_nxt_5_25_port);
   regs_reg_5_25_inst : DFF_X1 port map( D => N880, CK => clk, Q => 
                           regs_5_25_port, QN => n_1175);
   regs_nxt_reg_5_24_inst : DLH_X1 port map( G => n27505, D => n27417, Q => 
                           regs_nxt_5_24_port);
   regs_reg_5_24_inst : DFF_X1 port map( D => N879, CK => clk, Q => 
                           regs_5_24_port, QN => n_1176);
   regs_nxt_reg_5_23_inst : DLH_X1 port map( G => n27505, D => n27423, Q => 
                           regs_nxt_5_23_port);
   regs_reg_5_23_inst : DFF_X1 port map( D => N878, CK => clk, Q => 
                           regs_5_23_port, QN => n_1177);
   regs_nxt_reg_5_22_inst : DLH_X1 port map( G => n27505, D => n27429, Q => 
                           regs_nxt_5_22_port);
   regs_reg_5_22_inst : DFF_X1 port map( D => N877, CK => clk, Q => 
                           regs_5_22_port, QN => n_1178);
   regs_nxt_reg_5_21_inst : DLH_X1 port map( G => n27503, D => n27435, Q => 
                           regs_nxt_5_21_port);
   regs_reg_5_21_inst : DFF_X1 port map( D => N876, CK => clk, Q => 
                           regs_5_21_port, QN => n_1179);
   regs_nxt_reg_5_20_inst : DLH_X1 port map( G => n27503, D => n27285, Q => 
                           regs_nxt_5_20_port);
   regs_reg_5_20_inst : DFF_X1 port map( D => N875, CK => clk, Q => 
                           regs_5_20_port, QN => n_1180);
   regs_nxt_reg_5_19_inst : DLH_X1 port map( G => n27503, D => n27291, Q => 
                           regs_nxt_5_19_port);
   regs_reg_5_19_inst : DFF_X1 port map( D => N874, CK => clk, Q => 
                           regs_5_19_port, QN => n_1181);
   regs_nxt_reg_5_18_inst : DLH_X1 port map( G => n27505, D => n27297, Q => 
                           regs_nxt_5_18_port);
   regs_reg_5_18_inst : DFF_X1 port map( D => N873, CK => clk, Q => 
                           regs_5_18_port, QN => n_1182);
   regs_nxt_reg_5_17_inst : DLH_X1 port map( G => n27503, D => n27303, Q => 
                           regs_nxt_5_17_port);
   regs_reg_5_17_inst : DFF_X1 port map( D => N872, CK => clk, Q => 
                           regs_5_17_port, QN => n_1183);
   regs_nxt_reg_5_16_inst : DLH_X1 port map( G => n27505, D => n27309, Q => 
                           regs_nxt_5_16_port);
   regs_reg_5_16_inst : DFF_X1 port map( D => N871, CK => clk, Q => 
                           regs_5_16_port, QN => n_1184);
   regs_nxt_reg_5_15_inst : DLH_X1 port map( G => n27503, D => n27315, Q => 
                           regs_nxt_5_15_port);
   regs_reg_5_15_inst : DFF_X1 port map( D => N870, CK => clk, Q => 
                           regs_5_15_port, QN => n_1185);
   regs_nxt_reg_5_14_inst : DLH_X1 port map( G => n27505, D => n27321, Q => 
                           regs_nxt_5_14_port);
   regs_reg_5_14_inst : DFF_X1 port map( D => N869, CK => clk, Q => 
                           regs_5_14_port, QN => n_1186);
   regs_nxt_reg_5_13_inst : DLH_X1 port map( G => n27505, D => n27327, Q => 
                           regs_nxt_5_13_port);
   regs_reg_5_13_inst : DFF_X1 port map( D => N868, CK => clk, Q => 
                           regs_5_13_port, QN => n_1187);
   regs_nxt_reg_5_12_inst : DLH_X1 port map( G => n27505, D => n27333, Q => 
                           regs_nxt_5_12_port);
   regs_reg_5_12_inst : DFF_X1 port map( D => N867, CK => clk, Q => 
                           regs_5_12_port, QN => n_1188);
   regs_nxt_reg_5_11_inst : DLH_X1 port map( G => n27503, D => n27339, Q => 
                           regs_nxt_5_11_port);
   regs_reg_5_11_inst : DFF_X1 port map( D => N866, CK => clk, Q => 
                           regs_5_11_port, QN => n_1189);
   regs_nxt_reg_5_10_inst : DLH_X1 port map( G => n27503, D => n27345, Q => 
                           regs_nxt_5_10_port);
   regs_reg_5_10_inst : DFF_X1 port map( D => N865, CK => clk, Q => 
                           regs_5_10_port, QN => n_1190);
   regs_nxt_reg_5_9_inst : DLH_X1 port map( G => n27504, D => n27351, Q => 
                           regs_nxt_5_9_port);
   regs_reg_5_9_inst : DFF_X1 port map( D => N864, CK => clk, Q => 
                           regs_5_9_port, QN => n_1191);
   regs_nxt_reg_5_8_inst : DLH_X1 port map( G => n27504, D => n27357, Q => 
                           regs_nxt_5_8_port);
   regs_reg_5_8_inst : DFF_X1 port map( D => N863, CK => clk, Q => 
                           regs_5_8_port, QN => n_1192);
   regs_nxt_reg_5_7_inst : DLH_X1 port map( G => n27504, D => n27363, Q => 
                           regs_nxt_5_7_port);
   regs_reg_5_7_inst : DFF_X1 port map( D => N862, CK => clk, Q => 
                           regs_5_7_port, QN => n_1193);
   regs_nxt_reg_5_6_inst : DLH_X1 port map( G => n27504, D => n27369, Q => 
                           regs_nxt_5_6_port);
   regs_reg_5_6_inst : DFF_X1 port map( D => N861, CK => clk, Q => 
                           regs_5_6_port, QN => n_1194);
   regs_nxt_reg_5_5_inst : DLH_X1 port map( G => n27504, D => n27279, Q => 
                           regs_nxt_5_5_port);
   regs_reg_5_5_inst : DFF_X1 port map( D => N860, CK => clk, Q => 
                           regs_5_5_port, QN => n_1195);
   regs_nxt_reg_5_4_inst : DLH_X1 port map( G => n27504, D => n27441, Q => 
                           regs_nxt_5_4_port);
   regs_reg_5_4_inst : DFF_X1 port map( D => N859, CK => clk, Q => 
                           regs_5_4_port, QN => n_1196);
   regs_nxt_reg_5_3_inst : DLH_X1 port map( G => n27505, D => n27447, Q => 
                           regs_nxt_5_3_port);
   regs_reg_5_3_inst : DFF_X1 port map( D => N858, CK => clk, Q => 
                           regs_5_3_port, QN => n_1197);
   regs_nxt_reg_5_2_inst : DLH_X1 port map( G => n27504, D => n27453, Q => 
                           regs_nxt_5_2_port);
   regs_reg_5_2_inst : DFF_X1 port map( D => N857, CK => clk, Q => 
                           regs_5_2_port, QN => n_1198);
   regs_nxt_reg_5_1_inst : DLH_X1 port map( G => n27503, D => n27459, Q => 
                           regs_nxt_5_1_port);
   regs_reg_5_1_inst : DFF_X1 port map( D => N856, CK => clk, Q => 
                           regs_5_1_port, QN => n_1199);
   regs_nxt_reg_5_0_inst : DLH_X1 port map( G => n27504, D => n27465, Q => 
                           regs_nxt_5_0_port);
   regs_reg_5_0_inst : DFF_X1 port map( D => N855, CK => clk, Q => 
                           regs_5_0_port, QN => n_1200);
   regs_nxt_reg_6_31_inst : DLH_X1 port map( G => n27511, D => n27372, Q => 
                           regs_nxt_6_31_port);
   regs_reg_6_31_inst : DFF_X1 port map( D => N854, CK => clk, Q => n26425, QN 
                           => n2218);
   regs_nxt_reg_6_30_inst : DLH_X1 port map( G => n27511, D => n27378, Q => 
                           regs_nxt_6_30_port);
   regs_reg_6_30_inst : DFF_X1 port map( D => N853, CK => clk, Q => n26424, QN 
                           => n2211);
   regs_nxt_reg_6_29_inst : DLH_X1 port map( G => n27510, D => n27384, Q => 
                           regs_nxt_6_29_port);
   regs_reg_6_29_inst : DFF_X1 port map( D => N852, CK => clk, Q => n26423, QN 
                           => n2204);
   regs_nxt_reg_6_28_inst : DLH_X1 port map( G => n27510, D => n27390, Q => 
                           regs_nxt_6_28_port);
   regs_reg_6_28_inst : DFF_X1 port map( D => N851, CK => clk, Q => n26422, QN 
                           => n2197);
   regs_nxt_reg_6_27_inst : DLH_X1 port map( G => n27513, D => n27396, Q => 
                           regs_nxt_6_27_port);
   regs_reg_6_27_inst : DFF_X1 port map( D => N850, CK => clk, Q => n26421, QN 
                           => n2190);
   regs_nxt_reg_6_26_inst : DLH_X1 port map( G => n27512, D => n27402, Q => 
                           regs_nxt_6_26_port);
   regs_reg_6_26_inst : DFF_X1 port map( D => N849, CK => clk, Q => n26420, QN 
                           => n2183);
   regs_nxt_reg_6_25_inst : DLH_X1 port map( G => n27513, D => n27408, Q => 
                           regs_nxt_6_25_port);
   regs_reg_6_25_inst : DFF_X1 port map( D => N848, CK => clk, Q => n26419, QN 
                           => n2176);
   regs_nxt_reg_6_24_inst : DLH_X1 port map( G => n27512, D => n27414, Q => 
                           regs_nxt_6_24_port);
   regs_reg_6_24_inst : DFF_X1 port map( D => N847, CK => clk, Q => n26418, QN 
                           => n2169);
   regs_nxt_reg_6_23_inst : DLH_X1 port map( G => n27512, D => n27420, Q => 
                           regs_nxt_6_23_port);
   regs_reg_6_23_inst : DFF_X1 port map( D => N846, CK => clk, Q => n26417, QN 
                           => n2162);
   regs_nxt_reg_6_22_inst : DLH_X1 port map( G => n27512, D => n27426, Q => 
                           regs_nxt_6_22_port);
   regs_reg_6_22_inst : DFF_X1 port map( D => N845, CK => clk, Q => n26416, QN 
                           => n2155);
   regs_nxt_reg_6_21_inst : DLH_X1 port map( G => n27510, D => n27432, Q => 
                           regs_nxt_6_21_port);
   regs_reg_6_21_inst : DFF_X1 port map( D => N844, CK => clk, Q => n26415, QN 
                           => n2148);
   regs_nxt_reg_6_20_inst : DLH_X1 port map( G => n27510, D => n27282, Q => 
                           regs_nxt_6_20_port);
   regs_reg_6_20_inst : DFF_X1 port map( D => N843, CK => clk, Q => n26414, QN 
                           => n2141);
   regs_nxt_reg_6_19_inst : DLH_X1 port map( G => n27510, D => n27288, Q => 
                           regs_nxt_6_19_port);
   regs_reg_6_19_inst : DFF_X1 port map( D => N842, CK => clk, Q => n25485, QN 
                           => n_1201);
   regs_nxt_reg_6_18_inst : DLH_X1 port map( G => n27512, D => n27294, Q => 
                           regs_nxt_6_18_port);
   regs_reg_6_18_inst : DFF_X1 port map( D => N841, CK => clk, Q => n25484, QN 
                           => n_1202);
   regs_nxt_reg_6_17_inst : DLH_X1 port map( G => n27510, D => n27300, Q => 
                           regs_nxt_6_17_port);
   regs_reg_6_17_inst : DFF_X1 port map( D => N840, CK => clk, Q => n25483, QN 
                           => n_1203);
   regs_nxt_reg_6_16_inst : DLH_X1 port map( G => n27512, D => n27306, Q => 
                           regs_nxt_6_16_port);
   regs_reg_6_16_inst : DFF_X1 port map( D => N839, CK => clk, Q => n25482, QN 
                           => n_1204);
   regs_nxt_reg_6_15_inst : DLH_X1 port map( G => n27510, D => n27312, Q => 
                           regs_nxt_6_15_port);
   regs_reg_6_15_inst : DFF_X1 port map( D => N838, CK => clk, Q => n25481, QN 
                           => n_1205);
   regs_nxt_reg_6_14_inst : DLH_X1 port map( G => n27512, D => n27318, Q => 
                           regs_nxt_6_14_port);
   regs_reg_6_14_inst : DFF_X1 port map( D => N837, CK => clk, Q => n25480, QN 
                           => n_1206);
   regs_nxt_reg_6_13_inst : DLH_X1 port map( G => n27512, D => n27324, Q => 
                           regs_nxt_6_13_port);
   regs_reg_6_13_inst : DFF_X1 port map( D => N836, CK => clk, Q => n25479, QN 
                           => n_1207);
   regs_nxt_reg_6_12_inst : DLH_X1 port map( G => n27512, D => n27330, Q => 
                           regs_nxt_6_12_port);
   regs_reg_6_12_inst : DFF_X1 port map( D => N835, CK => clk, Q => n25478, QN 
                           => n_1208);
   regs_nxt_reg_6_11_inst : DLH_X1 port map( G => n27510, D => n27336, Q => 
                           regs_nxt_6_11_port);
   regs_reg_6_11_inst : DFF_X1 port map( D => N834, CK => clk, Q => n25477, QN 
                           => n_1209);
   regs_nxt_reg_6_10_inst : DLH_X1 port map( G => n27510, D => n27342, Q => 
                           regs_nxt_6_10_port);
   regs_reg_6_10_inst : DFF_X1 port map( D => N833, CK => clk, Q => n25476, QN 
                           => n_1210);
   regs_nxt_reg_6_9_inst : DLH_X1 port map( G => n27511, D => n27348, Q => 
                           regs_nxt_6_9_port);
   regs_reg_6_9_inst : DFF_X1 port map( D => N832, CK => clk, Q => n25475, QN 
                           => n_1211);
   regs_nxt_reg_6_8_inst : DLH_X1 port map( G => n27511, D => n27354, Q => 
                           regs_nxt_6_8_port);
   regs_reg_6_8_inst : DFF_X1 port map( D => N831, CK => clk, Q => n25474, QN 
                           => n_1212);
   regs_nxt_reg_6_7_inst : DLH_X1 port map( G => n27511, D => n27360, Q => 
                           regs_nxt_6_7_port);
   regs_reg_6_7_inst : DFF_X1 port map( D => N830, CK => clk, Q => n25473, QN 
                           => n_1213);
   regs_nxt_reg_6_6_inst : DLH_X1 port map( G => n27511, D => n27366, Q => 
                           regs_nxt_6_6_port);
   regs_reg_6_6_inst : DFF_X1 port map( D => N829, CK => clk, Q => n25472, QN 
                           => n_1214);
   regs_nxt_reg_6_5_inst : DLH_X1 port map( G => n27511, D => n27276, Q => 
                           regs_nxt_6_5_port);
   regs_reg_6_5_inst : DFF_X1 port map( D => N828, CK => clk, Q => n25471, QN 
                           => n_1215);
   regs_nxt_reg_6_4_inst : DLH_X1 port map( G => n27511, D => n27438, Q => 
                           regs_nxt_6_4_port);
   regs_reg_6_4_inst : DFF_X1 port map( D => N827, CK => clk, Q => n25470, QN 
                           => n_1216);
   regs_nxt_reg_6_3_inst : DLH_X1 port map( G => n27512, D => n27444, Q => 
                           regs_nxt_6_3_port);
   regs_reg_6_3_inst : DFF_X1 port map( D => N826, CK => clk, Q => n25469, QN 
                           => n_1217);
   regs_nxt_reg_6_2_inst : DLH_X1 port map( G => n27511, D => n27450, Q => 
                           regs_nxt_6_2_port);
   regs_reg_6_2_inst : DFF_X1 port map( D => N825, CK => clk, Q => n25468, QN 
                           => n_1218);
   regs_nxt_reg_6_1_inst : DLH_X1 port map( G => n27510, D => n27456, Q => 
                           regs_nxt_6_1_port);
   regs_reg_6_1_inst : DFF_X1 port map( D => N824, CK => clk, Q => n25467, QN 
                           => n_1219);
   regs_nxt_reg_6_0_inst : DLH_X1 port map( G => n27511, D => n27462, Q => 
                           regs_nxt_6_0_port);
   regs_reg_6_0_inst : DFF_X1 port map( D => N823, CK => clk, Q => n25466, QN 
                           => n_1220);
   regs_nxt_reg_7_31_inst : DLH_X1 port map( G => n27518, D => n27372, Q => 
                           regs_nxt_7_31_port);
   regs_reg_7_31_inst : DFF_X1 port map( D => N822, CK => clk, Q => 
                           regs_7_31_port, QN => n_1221);
   regs_nxt_reg_7_30_inst : DLH_X1 port map( G => n27518, D => n27378, Q => 
                           regs_nxt_7_30_port);
   regs_reg_7_30_inst : DFF_X1 port map( D => N821, CK => clk, Q => 
                           regs_7_30_port, QN => n_1222);
   regs_nxt_reg_7_29_inst : DLH_X1 port map( G => n27517, D => n27384, Q => 
                           regs_nxt_7_29_port);
   regs_reg_7_29_inst : DFF_X1 port map( D => N820, CK => clk, Q => 
                           regs_7_29_port, QN => n_1223);
   regs_nxt_reg_7_28_inst : DLH_X1 port map( G => n27517, D => n27390, Q => 
                           regs_nxt_7_28_port);
   regs_reg_7_28_inst : DFF_X1 port map( D => N819, CK => clk, Q => 
                           regs_7_28_port, QN => n_1224);
   regs_nxt_reg_7_27_inst : DLH_X1 port map( G => n27520, D => n27396, Q => 
                           regs_nxt_7_27_port);
   regs_reg_7_27_inst : DFF_X1 port map( D => N818, CK => clk, Q => 
                           regs_7_27_port, QN => n_1225);
   regs_nxt_reg_7_26_inst : DLH_X1 port map( G => n27519, D => n27402, Q => 
                           regs_nxt_7_26_port);
   regs_reg_7_26_inst : DFF_X1 port map( D => N817, CK => clk, Q => 
                           regs_7_26_port, QN => n_1226);
   regs_nxt_reg_7_25_inst : DLH_X1 port map( G => n27520, D => n27408, Q => 
                           regs_nxt_7_25_port);
   regs_reg_7_25_inst : DFF_X1 port map( D => N816, CK => clk, Q => 
                           regs_7_25_port, QN => n_1227);
   regs_nxt_reg_7_24_inst : DLH_X1 port map( G => n27519, D => n27414, Q => 
                           regs_nxt_7_24_port);
   regs_reg_7_24_inst : DFF_X1 port map( D => N815, CK => clk, Q => 
                           regs_7_24_port, QN => n_1228);
   regs_nxt_reg_7_23_inst : DLH_X1 port map( G => n27519, D => n27420, Q => 
                           regs_nxt_7_23_port);
   regs_reg_7_23_inst : DFF_X1 port map( D => N814, CK => clk, Q => 
                           regs_7_23_port, QN => n_1229);
   regs_nxt_reg_7_22_inst : DLH_X1 port map( G => n27519, D => n27426, Q => 
                           regs_nxt_7_22_port);
   regs_reg_7_22_inst : DFF_X1 port map( D => N813, CK => clk, Q => 
                           regs_7_22_port, QN => n_1230);
   regs_nxt_reg_7_21_inst : DLH_X1 port map( G => n27517, D => n27432, Q => 
                           regs_nxt_7_21_port);
   regs_reg_7_21_inst : DFF_X1 port map( D => N812, CK => clk, Q => 
                           regs_7_21_port, QN => n_1231);
   regs_nxt_reg_7_20_inst : DLH_X1 port map( G => n27517, D => n27282, Q => 
                           regs_nxt_7_20_port);
   regs_reg_7_20_inst : DFF_X1 port map( D => N811, CK => clk, Q => 
                           regs_7_20_port, QN => n_1232);
   regs_nxt_reg_7_19_inst : DLH_X1 port map( G => n27517, D => n27288, Q => 
                           regs_nxt_7_19_port);
   regs_reg_7_19_inst : DFF_X1 port map( D => N810, CK => clk, Q => 
                           regs_7_19_port, QN => n_1233);
   regs_nxt_reg_7_18_inst : DLH_X1 port map( G => n27519, D => n27294, Q => 
                           regs_nxt_7_18_port);
   regs_reg_7_18_inst : DFF_X1 port map( D => N809, CK => clk, Q => 
                           regs_7_18_port, QN => n_1234);
   regs_nxt_reg_7_17_inst : DLH_X1 port map( G => n27517, D => n27300, Q => 
                           regs_nxt_7_17_port);
   regs_reg_7_17_inst : DFF_X1 port map( D => N808, CK => clk, Q => 
                           regs_7_17_port, QN => n_1235);
   regs_nxt_reg_7_16_inst : DLH_X1 port map( G => n27519, D => n27306, Q => 
                           regs_nxt_7_16_port);
   regs_reg_7_16_inst : DFF_X1 port map( D => N807, CK => clk, Q => 
                           regs_7_16_port, QN => n_1236);
   regs_nxt_reg_7_15_inst : DLH_X1 port map( G => n27517, D => n27312, Q => 
                           regs_nxt_7_15_port);
   regs_reg_7_15_inst : DFF_X1 port map( D => N806, CK => clk, Q => 
                           regs_7_15_port, QN => n_1237);
   regs_nxt_reg_7_14_inst : DLH_X1 port map( G => n27519, D => n27318, Q => 
                           regs_nxt_7_14_port);
   regs_reg_7_14_inst : DFF_X1 port map( D => N805, CK => clk, Q => 
                           regs_7_14_port, QN => n_1238);
   regs_nxt_reg_7_13_inst : DLH_X1 port map( G => n27519, D => n27324, Q => 
                           regs_nxt_7_13_port);
   regs_reg_7_13_inst : DFF_X1 port map( D => N804, CK => clk, Q => 
                           regs_7_13_port, QN => n_1239);
   regs_nxt_reg_7_12_inst : DLH_X1 port map( G => n27519, D => n27330, Q => 
                           regs_nxt_7_12_port);
   regs_reg_7_12_inst : DFF_X1 port map( D => N803, CK => clk, Q => 
                           regs_7_12_port, QN => n_1240);
   regs_nxt_reg_7_11_inst : DLH_X1 port map( G => n27517, D => n27336, Q => 
                           regs_nxt_7_11_port);
   regs_reg_7_11_inst : DFF_X1 port map( D => N802, CK => clk, Q => 
                           regs_7_11_port, QN => n_1241);
   regs_nxt_reg_7_10_inst : DLH_X1 port map( G => n27517, D => n27342, Q => 
                           regs_nxt_7_10_port);
   regs_reg_7_10_inst : DFF_X1 port map( D => N801, CK => clk, Q => 
                           regs_7_10_port, QN => n_1242);
   regs_nxt_reg_7_9_inst : DLH_X1 port map( G => n27518, D => n27348, Q => 
                           regs_nxt_7_9_port);
   regs_reg_7_9_inst : DFF_X1 port map( D => N800, CK => clk, Q => 
                           regs_7_9_port, QN => n_1243);
   regs_nxt_reg_7_8_inst : DLH_X1 port map( G => n27518, D => n27354, Q => 
                           regs_nxt_7_8_port);
   regs_reg_7_8_inst : DFF_X1 port map( D => N799, CK => clk, Q => 
                           regs_7_8_port, QN => n_1244);
   regs_nxt_reg_7_7_inst : DLH_X1 port map( G => n27518, D => n27360, Q => 
                           regs_nxt_7_7_port);
   regs_reg_7_7_inst : DFF_X1 port map( D => N798, CK => clk, Q => 
                           regs_7_7_port, QN => n_1245);
   regs_nxt_reg_7_6_inst : DLH_X1 port map( G => n27518, D => n27366, Q => 
                           regs_nxt_7_6_port);
   regs_reg_7_6_inst : DFF_X1 port map( D => N797, CK => clk, Q => 
                           regs_7_6_port, QN => n_1246);
   regs_nxt_reg_7_5_inst : DLH_X1 port map( G => n27518, D => n27276, Q => 
                           regs_nxt_7_5_port);
   regs_reg_7_5_inst : DFF_X1 port map( D => N796, CK => clk, Q => 
                           regs_7_5_port, QN => n_1247);
   regs_nxt_reg_7_4_inst : DLH_X1 port map( G => n27518, D => n27438, Q => 
                           regs_nxt_7_4_port);
   regs_reg_7_4_inst : DFF_X1 port map( D => N795, CK => clk, Q => 
                           regs_7_4_port, QN => n_1248);
   regs_nxt_reg_7_3_inst : DLH_X1 port map( G => n27519, D => n27444, Q => 
                           regs_nxt_7_3_port);
   regs_reg_7_3_inst : DFF_X1 port map( D => N794, CK => clk, Q => 
                           regs_7_3_port, QN => n_1249);
   regs_nxt_reg_7_2_inst : DLH_X1 port map( G => n27518, D => n27450, Q => 
                           regs_nxt_7_2_port);
   regs_reg_7_2_inst : DFF_X1 port map( D => N793, CK => clk, Q => 
                           regs_7_2_port, QN => n_1250);
   regs_nxt_reg_7_1_inst : DLH_X1 port map( G => n27517, D => n27456, Q => 
                           regs_nxt_7_1_port);
   regs_reg_7_1_inst : DFF_X1 port map( D => N792, CK => clk, Q => 
                           regs_7_1_port, QN => n_1251);
   regs_nxt_reg_7_0_inst : DLH_X1 port map( G => n27518, D => n27462, Q => 
                           regs_nxt_7_0_port);
   regs_reg_7_0_inst : DFF_X1 port map( D => N791, CK => clk, Q => 
                           regs_7_0_port, QN => n_1252);
   regs_nxt_reg_8_31_inst : DLH_X1 port map( G => n27525, D => n27372, Q => 
                           regs_nxt_8_31_port);
   regs_reg_8_31_inst : DFF_X1 port map( D => N790, CK => clk, Q => n_1253, QN 
                           => n26631);
   regs_nxt_reg_8_30_inst : DLH_X1 port map( G => n27525, D => n27380, Q => 
                           regs_nxt_8_30_port);
   regs_reg_8_30_inst : DFF_X1 port map( D => N789, CK => clk, Q => n_1254, QN 
                           => n26630);
   regs_nxt_reg_8_29_inst : DLH_X1 port map( G => n27524, D => n27384, Q => 
                           regs_nxt_8_29_port);
   regs_reg_8_29_inst : DFF_X1 port map( D => N788, CK => clk, Q => n_1255, QN 
                           => n26629);
   regs_nxt_reg_8_28_inst : DLH_X1 port map( G => n27524, D => n27392, Q => 
                           regs_nxt_8_28_port);
   regs_reg_8_28_inst : DFF_X1 port map( D => N787, CK => clk, Q => n_1256, QN 
                           => n26628);
   regs_nxt_reg_8_27_inst : DLH_X1 port map( G => n27524, D => n27396, Q => 
                           regs_nxt_8_27_port);
   regs_reg_8_27_inst : DFF_X1 port map( D => N786, CK => clk, Q => n_1257, QN 
                           => n26627);
   regs_nxt_reg_8_26_inst : DLH_X1 port map( G => n27526, D => n27404, Q => 
                           regs_nxt_8_26_port);
   regs_reg_8_26_inst : DFF_X1 port map( D => N785, CK => clk, Q => n_1258, QN 
                           => n26626);
   regs_nxt_reg_8_25_inst : DLH_X1 port map( G => n27527, D => n27408, Q => 
                           regs_nxt_8_25_port);
   regs_reg_8_25_inst : DFF_X1 port map( D => N784, CK => clk, Q => n_1259, QN 
                           => n26625);
   regs_nxt_reg_8_24_inst : DLH_X1 port map( G => n27526, D => n27416, Q => 
                           regs_nxt_8_24_port);
   regs_reg_8_24_inst : DFF_X1 port map( D => N783, CK => clk, Q => n_1260, QN 
                           => n26624);
   regs_nxt_reg_8_23_inst : DLH_X1 port map( G => n27527, D => n27420, Q => 
                           regs_nxt_8_23_port);
   regs_reg_8_23_inst : DFF_X1 port map( D => N782, CK => clk, Q => n_1261, QN 
                           => n26623);
   regs_nxt_reg_8_22_inst : DLH_X1 port map( G => n27526, D => n27428, Q => 
                           regs_nxt_8_22_port);
   regs_reg_8_22_inst : DFF_X1 port map( D => N781, CK => clk, Q => n_1262, QN 
                           => n26622);
   regs_nxt_reg_8_21_inst : DLH_X1 port map( G => n27526, D => n27432, Q => 
                           regs_nxt_8_21_port);
   regs_reg_8_21_inst : DFF_X1 port map( D => N780, CK => clk, Q => n_1263, QN 
                           => n26621);
   regs_nxt_reg_8_20_inst : DLH_X1 port map( G => n27524, D => n27284, Q => 
                           regs_nxt_8_20_port);
   regs_reg_8_20_inst : DFF_X1 port map( D => N779, CK => clk, Q => n_1264, QN 
                           => n26620);
   regs_nxt_reg_8_19_inst : DLH_X1 port map( G => n27524, D => n27288, Q => 
                           regs_nxt_8_19_port);
   regs_reg_8_19_inst : DFF_X1 port map( D => N778, CK => clk, Q => n_1265, QN 
                           => n26619);
   regs_nxt_reg_8_18_inst : DLH_X1 port map( G => n27526, D => n27296, Q => 
                           regs_nxt_8_18_port);
   regs_reg_8_18_inst : DFF_X1 port map( D => N777, CK => clk, Q => n_1266, QN 
                           => n26618);
   regs_nxt_reg_8_17_inst : DLH_X1 port map( G => n27524, D => n27300, Q => 
                           regs_nxt_8_17_port);
   regs_reg_8_17_inst : DFF_X1 port map( D => N776, CK => clk, Q => n_1267, QN 
                           => n26617);
   regs_nxt_reg_8_16_inst : DLH_X1 port map( G => n27526, D => n27308, Q => 
                           regs_nxt_8_16_port);
   regs_reg_8_16_inst : DFF_X1 port map( D => N775, CK => clk, Q => n_1268, QN 
                           => n26616);
   regs_nxt_reg_8_15_inst : DLH_X1 port map( G => n27524, D => n27312, Q => 
                           regs_nxt_8_15_port);
   regs_reg_8_15_inst : DFF_X1 port map( D => N774, CK => clk, Q => n_1269, QN 
                           => n26615);
   regs_nxt_reg_8_14_inst : DLH_X1 port map( G => n27526, D => n27320, Q => 
                           regs_nxt_8_14_port);
   regs_reg_8_14_inst : DFF_X1 port map( D => N773, CK => clk, Q => n_1270, QN 
                           => n26614);
   regs_nxt_reg_8_13_inst : DLH_X1 port map( G => n27526, D => n27324, Q => 
                           regs_nxt_8_13_port);
   regs_reg_8_13_inst : DFF_X1 port map( D => N772, CK => clk, Q => n_1271, QN 
                           => n26613);
   regs_nxt_reg_8_12_inst : DLH_X1 port map( G => n27526, D => n27332, Q => 
                           regs_nxt_8_12_port);
   regs_reg_8_12_inst : DFF_X1 port map( D => N771, CK => clk, Q => n_1272, QN 
                           => n26612);
   regs_nxt_reg_8_11_inst : DLH_X1 port map( G => n27524, D => n27336, Q => 
                           regs_nxt_8_11_port);
   regs_reg_8_11_inst : DFF_X1 port map( D => N770, CK => clk, Q => n_1273, QN 
                           => n26611);
   regs_nxt_reg_8_10_inst : DLH_X1 port map( G => n27524, D => n27344, Q => 
                           regs_nxt_8_10_port);
   regs_reg_8_10_inst : DFF_X1 port map( D => N769, CK => clk, Q => n_1274, QN 
                           => n26610);
   regs_nxt_reg_8_9_inst : DLH_X1 port map( G => n27525, D => n27348, Q => 
                           regs_nxt_8_9_port);
   regs_reg_8_9_inst : DFF_X1 port map( D => N768, CK => clk, Q => n_1275, QN 
                           => n26609);
   regs_nxt_reg_8_8_inst : DLH_X1 port map( G => n27525, D => n27356, Q => 
                           regs_nxt_8_8_port);
   regs_reg_8_8_inst : DFF_X1 port map( D => N767, CK => clk, Q => n_1276, QN 
                           => n26608);
   regs_nxt_reg_8_7_inst : DLH_X1 port map( G => n27525, D => n27360, Q => 
                           regs_nxt_8_7_port);
   regs_reg_8_7_inst : DFF_X1 port map( D => N766, CK => clk, Q => n_1277, QN 
                           => n26607);
   regs_nxt_reg_8_6_inst : DLH_X1 port map( G => n27525, D => n27368, Q => 
                           regs_nxt_8_6_port);
   regs_reg_8_6_inst : DFF_X1 port map( D => N765, CK => clk, Q => n_1278, QN 
                           => n26606);
   regs_nxt_reg_8_5_inst : DLH_X1 port map( G => n27525, D => n27278, Q => 
                           regs_nxt_8_5_port);
   regs_reg_8_5_inst : DFF_X1 port map( D => N764, CK => clk, Q => n_1279, QN 
                           => n26605);
   regs_nxt_reg_8_4_inst : DLH_X1 port map( G => n27525, D => n27440, Q => 
                           regs_nxt_8_4_port);
   regs_reg_8_4_inst : DFF_X1 port map( D => N763, CK => clk, Q => n_1280, QN 
                           => n26604);
   regs_nxt_reg_8_3_inst : DLH_X1 port map( G => n27526, D => n27444, Q => 
                           regs_nxt_8_3_port);
   regs_reg_8_3_inst : DFF_X1 port map( D => N762, CK => clk, Q => n_1281, QN 
                           => n26603);
   regs_nxt_reg_8_2_inst : DLH_X1 port map( G => n27525, D => n27450, Q => 
                           regs_nxt_8_2_port);
   regs_reg_8_2_inst : DFF_X1 port map( D => N761, CK => clk, Q => n_1282, QN 
                           => n26602);
   regs_nxt_reg_8_1_inst : DLH_X1 port map( G => n27524, D => n27456, Q => 
                           regs_nxt_8_1_port);
   regs_reg_8_1_inst : DFF_X1 port map( D => N760, CK => clk, Q => n_1283, QN 
                           => n26601);
   regs_nxt_reg_8_0_inst : DLH_X1 port map( G => n27525, D => n27464, Q => 
                           regs_nxt_8_0_port);
   regs_reg_8_0_inst : DFF_X1 port map( D => N759, CK => clk, Q => n_1284, QN 
                           => n26600);
   regs_nxt_reg_9_31_inst : DLH_X1 port map( G => n27532, D => n27374, Q => 
                           regs_nxt_9_31_port);
   regs_reg_9_31_inst : DFF_X1 port map( D => N758, CK => clk, Q => n_1285, QN 
                           => n26663);
   regs_nxt_reg_9_30_inst : DLH_X1 port map( G => n27532, D => n27378, Q => 
                           regs_nxt_9_30_port);
   regs_reg_9_30_inst : DFF_X1 port map( D => N757, CK => clk, Q => n_1286, QN 
                           => n26662);
   regs_nxt_reg_9_29_inst : DLH_X1 port map( G => n27531, D => n27386, Q => 
                           regs_nxt_9_29_port);
   regs_reg_9_29_inst : DFF_X1 port map( D => N756, CK => clk, Q => n_1287, QN 
                           => n26661);
   regs_nxt_reg_9_28_inst : DLH_X1 port map( G => n27531, D => n27390, Q => 
                           regs_nxt_9_28_port);
   regs_reg_9_28_inst : DFF_X1 port map( D => N755, CK => clk, Q => n_1288, QN 
                           => n26660);
   regs_nxt_reg_9_27_inst : DLH_X1 port map( G => n27534, D => n27398, Q => 
                           regs_nxt_9_27_port);
   regs_reg_9_27_inst : DFF_X1 port map( D => N754, CK => clk, Q => n_1289, QN 
                           => n26659);
   regs_nxt_reg_9_26_inst : DLH_X1 port map( G => n27533, D => n27402, Q => 
                           regs_nxt_9_26_port);
   regs_reg_9_26_inst : DFF_X1 port map( D => N753, CK => clk, Q => n_1290, QN 
                           => n26658);
   regs_nxt_reg_9_25_inst : DLH_X1 port map( G => n27534, D => n27410, Q => 
                           regs_nxt_9_25_port);
   regs_reg_9_25_inst : DFF_X1 port map( D => N752, CK => clk, Q => n_1291, QN 
                           => n26657);
   regs_nxt_reg_9_24_inst : DLH_X1 port map( G => n27533, D => n27414, Q => 
                           regs_nxt_9_24_port);
   regs_reg_9_24_inst : DFF_X1 port map( D => N751, CK => clk, Q => n_1292, QN 
                           => n26656);
   regs_nxt_reg_9_23_inst : DLH_X1 port map( G => n27533, D => n27422, Q => 
                           regs_nxt_9_23_port);
   regs_reg_9_23_inst : DFF_X1 port map( D => N750, CK => clk, Q => n_1293, QN 
                           => n26655);
   regs_nxt_reg_9_22_inst : DLH_X1 port map( G => n27533, D => n27426, Q => 
                           regs_nxt_9_22_port);
   regs_reg_9_22_inst : DFF_X1 port map( D => N749, CK => clk, Q => n_1294, QN 
                           => n26654);
   regs_nxt_reg_9_21_inst : DLH_X1 port map( G => n27531, D => n27434, Q => 
                           regs_nxt_9_21_port);
   regs_reg_9_21_inst : DFF_X1 port map( D => N748, CK => clk, Q => n_1295, QN 
                           => n26653);
   regs_nxt_reg_9_20_inst : DLH_X1 port map( G => n27531, D => n27282, Q => 
                           regs_nxt_9_20_port);
   regs_reg_9_20_inst : DFF_X1 port map( D => N747, CK => clk, Q => n_1296, QN 
                           => n26652);
   regs_nxt_reg_9_19_inst : DLH_X1 port map( G => n27531, D => n27290, Q => 
                           regs_nxt_9_19_port);
   regs_reg_9_19_inst : DFF_X1 port map( D => N746, CK => clk, Q => n_1297, QN 
                           => n26651);
   regs_nxt_reg_9_18_inst : DLH_X1 port map( G => n27533, D => n27294, Q => 
                           regs_nxt_9_18_port);
   regs_reg_9_18_inst : DFF_X1 port map( D => N745, CK => clk, Q => n_1298, QN 
                           => n26650);
   regs_nxt_reg_9_17_inst : DLH_X1 port map( G => n27531, D => n27302, Q => 
                           regs_nxt_9_17_port);
   regs_reg_9_17_inst : DFF_X1 port map( D => N744, CK => clk, Q => n_1299, QN 
                           => n26649);
   regs_nxt_reg_9_16_inst : DLH_X1 port map( G => n27533, D => n27306, Q => 
                           regs_nxt_9_16_port);
   regs_reg_9_16_inst : DFF_X1 port map( D => N743, CK => clk, Q => n_1300, QN 
                           => n26648);
   regs_nxt_reg_9_15_inst : DLH_X1 port map( G => n27531, D => n27314, Q => 
                           regs_nxt_9_15_port);
   regs_reg_9_15_inst : DFF_X1 port map( D => N742, CK => clk, Q => n_1301, QN 
                           => n26647);
   regs_nxt_reg_9_14_inst : DLH_X1 port map( G => n27533, D => n27318, Q => 
                           regs_nxt_9_14_port);
   regs_reg_9_14_inst : DFF_X1 port map( D => N741, CK => clk, Q => n_1302, QN 
                           => n26646);
   regs_nxt_reg_9_13_inst : DLH_X1 port map( G => n27533, D => n27326, Q => 
                           regs_nxt_9_13_port);
   regs_reg_9_13_inst : DFF_X1 port map( D => N740, CK => clk, Q => n_1303, QN 
                           => n26645);
   regs_nxt_reg_9_12_inst : DLH_X1 port map( G => n27533, D => n27330, Q => 
                           regs_nxt_9_12_port);
   regs_reg_9_12_inst : DFF_X1 port map( D => N739, CK => clk, Q => n_1304, QN 
                           => n26644);
   regs_nxt_reg_9_11_inst : DLH_X1 port map( G => n27531, D => n27338, Q => 
                           regs_nxt_9_11_port);
   regs_reg_9_11_inst : DFF_X1 port map( D => N738, CK => clk, Q => n_1305, QN 
                           => n26643);
   regs_nxt_reg_9_10_inst : DLH_X1 port map( G => n27531, D => n27342, Q => 
                           regs_nxt_9_10_port);
   regs_reg_9_10_inst : DFF_X1 port map( D => N737, CK => clk, Q => n_1306, QN 
                           => n26642);
   regs_nxt_reg_9_9_inst : DLH_X1 port map( G => n27532, D => n27350, Q => 
                           regs_nxt_9_9_port);
   regs_reg_9_9_inst : DFF_X1 port map( D => N736, CK => clk, Q => n_1307, QN 
                           => n26641);
   regs_nxt_reg_9_8_inst : DLH_X1 port map( G => n27532, D => n27354, Q => 
                           regs_nxt_9_8_port);
   regs_reg_9_8_inst : DFF_X1 port map( D => N735, CK => clk, Q => n_1308, QN 
                           => n26640);
   regs_nxt_reg_9_7_inst : DLH_X1 port map( G => n27532, D => n27362, Q => 
                           regs_nxt_9_7_port);
   regs_reg_9_7_inst : DFF_X1 port map( D => N734, CK => clk, Q => n_1309, QN 
                           => n26639);
   regs_nxt_reg_9_6_inst : DLH_X1 port map( G => n27532, D => n27366, Q => 
                           regs_nxt_9_6_port);
   regs_reg_9_6_inst : DFF_X1 port map( D => N733, CK => clk, Q => n_1310, QN 
                           => n26638);
   regs_nxt_reg_9_5_inst : DLH_X1 port map( G => n27532, D => n27276, Q => 
                           regs_nxt_9_5_port);
   regs_reg_9_5_inst : DFF_X1 port map( D => N732, CK => clk, Q => n_1311, QN 
                           => n26637);
   regs_nxt_reg_9_4_inst : DLH_X1 port map( G => n27532, D => n27438, Q => 
                           regs_nxt_9_4_port);
   regs_reg_9_4_inst : DFF_X1 port map( D => N731, CK => clk, Q => n_1312, QN 
                           => n26636);
   regs_nxt_reg_9_3_inst : DLH_X1 port map( G => n27533, D => n27446, Q => 
                           regs_nxt_9_3_port);
   regs_reg_9_3_inst : DFF_X1 port map( D => N730, CK => clk, Q => n_1313, QN 
                           => n26635);
   regs_nxt_reg_9_2_inst : DLH_X1 port map( G => n27532, D => n27452, Q => 
                           regs_nxt_9_2_port);
   regs_reg_9_2_inst : DFF_X1 port map( D => N729, CK => clk, Q => n_1314, QN 
                           => n26634);
   regs_nxt_reg_9_1_inst : DLH_X1 port map( G => n27531, D => n27458, Q => 
                           regs_nxt_9_1_port);
   regs_reg_9_1_inst : DFF_X1 port map( D => N728, CK => clk, Q => n_1315, QN 
                           => n26633);
   regs_nxt_reg_9_0_inst : DLH_X1 port map( G => n27532, D => n27462, Q => 
                           regs_nxt_9_0_port);
   regs_reg_9_0_inst : DFF_X1 port map( D => N727, CK => clk, Q => n_1316, QN 
                           => n26632);
   regs_nxt_reg_10_31_inst : DLH_X1 port map( G => n27539, D => n27374, Q => 
                           regs_nxt_10_31_port);
   regs_reg_10_31_inst : DFF_X1 port map( D => N726, CK => clk, Q => n2217, QN 
                           => n26888);
   regs_nxt_reg_10_30_inst : DLH_X1 port map( G => n27539, D => n27380, Q => 
                           regs_nxt_10_30_port);
   regs_reg_10_30_inst : DFF_X1 port map( D => N725, CK => clk, Q => n2210, QN 
                           => n26886);
   regs_nxt_reg_10_29_inst : DLH_X1 port map( G => n27538, D => n27386, Q => 
                           regs_nxt_10_29_port);
   regs_reg_10_29_inst : DFF_X1 port map( D => N724, CK => clk, Q => n2203, QN 
                           => n26884);
   regs_nxt_reg_10_28_inst : DLH_X1 port map( G => n27538, D => n27392, Q => 
                           regs_nxt_10_28_port);
   regs_reg_10_28_inst : DFF_X1 port map( D => N723, CK => clk, Q => n2196, QN 
                           => n26882);
   regs_nxt_reg_10_27_inst : DLH_X1 port map( G => n27541, D => n27398, Q => 
                           regs_nxt_10_27_port);
   regs_reg_10_27_inst : DFF_X1 port map( D => N722, CK => clk, Q => n2189, QN 
                           => n26880);
   regs_nxt_reg_10_26_inst : DLH_X1 port map( G => n27540, D => n27404, Q => 
                           regs_nxt_10_26_port);
   regs_reg_10_26_inst : DFF_X1 port map( D => N721, CK => clk, Q => n2182, QN 
                           => n26878);
   regs_nxt_reg_10_25_inst : DLH_X1 port map( G => n27541, D => n27410, Q => 
                           regs_nxt_10_25_port);
   regs_reg_10_25_inst : DFF_X1 port map( D => N720, CK => clk, Q => n2175, QN 
                           => n26876);
   regs_nxt_reg_10_24_inst : DLH_X1 port map( G => n27540, D => n27416, Q => 
                           regs_nxt_10_24_port);
   regs_reg_10_24_inst : DFF_X1 port map( D => N719, CK => clk, Q => n2168, QN 
                           => n26874);
   regs_nxt_reg_10_23_inst : DLH_X1 port map( G => n27540, D => n27422, Q => 
                           regs_nxt_10_23_port);
   regs_reg_10_23_inst : DFF_X1 port map( D => N718, CK => clk, Q => n2161, QN 
                           => n26872);
   regs_nxt_reg_10_22_inst : DLH_X1 port map( G => n27540, D => n27428, Q => 
                           regs_nxt_10_22_port);
   regs_reg_10_22_inst : DFF_X1 port map( D => N717, CK => clk, Q => n2154, QN 
                           => n26870);
   regs_nxt_reg_10_21_inst : DLH_X1 port map( G => n27538, D => n27434, Q => 
                           regs_nxt_10_21_port);
   regs_reg_10_21_inst : DFF_X1 port map( D => N716, CK => clk, Q => n2147, QN 
                           => n26868);
   regs_nxt_reg_10_20_inst : DLH_X1 port map( G => n27538, D => n27284, Q => 
                           regs_nxt_10_20_port);
   regs_reg_10_20_inst : DFF_X1 port map( D => N715, CK => clk, Q => n2140, QN 
                           => n26866);
   regs_nxt_reg_10_19_inst : DLH_X1 port map( G => n27538, D => n27290, Q => 
                           regs_nxt_10_19_port);
   regs_reg_10_19_inst : DFF_X1 port map( D => N714, CK => clk, Q => n_1317, QN
                           => n25310);
   regs_nxt_reg_10_18_inst : DLH_X1 port map( G => n27540, D => n27296, Q => 
                           regs_nxt_10_18_port);
   regs_reg_10_18_inst : DFF_X1 port map( D => N713, CK => clk, Q => n_1318, QN
                           => n25309);
   regs_nxt_reg_10_17_inst : DLH_X1 port map( G => n27538, D => n27302, Q => 
                           regs_nxt_10_17_port);
   regs_reg_10_17_inst : DFF_X1 port map( D => N712, CK => clk, Q => n_1319, QN
                           => n25308);
   regs_nxt_reg_10_16_inst : DLH_X1 port map( G => n27540, D => n27308, Q => 
                           regs_nxt_10_16_port);
   regs_reg_10_16_inst : DFF_X1 port map( D => N711, CK => clk, Q => n_1320, QN
                           => n25307);
   regs_nxt_reg_10_15_inst : DLH_X1 port map( G => n27538, D => n27314, Q => 
                           regs_nxt_10_15_port);
   regs_reg_10_15_inst : DFF_X1 port map( D => N710, CK => clk, Q => n_1321, QN
                           => n25306);
   regs_nxt_reg_10_14_inst : DLH_X1 port map( G => n27540, D => n27320, Q => 
                           regs_nxt_10_14_port);
   regs_reg_10_14_inst : DFF_X1 port map( D => N709, CK => clk, Q => n_1322, QN
                           => n25305);
   regs_nxt_reg_10_13_inst : DLH_X1 port map( G => n27540, D => n27326, Q => 
                           regs_nxt_10_13_port);
   regs_reg_10_13_inst : DFF_X1 port map( D => N708, CK => clk, Q => n_1323, QN
                           => n25304);
   regs_nxt_reg_10_12_inst : DLH_X1 port map( G => n27540, D => n27332, Q => 
                           regs_nxt_10_12_port);
   regs_reg_10_12_inst : DFF_X1 port map( D => N707, CK => clk, Q => n_1324, QN
                           => n25303);
   regs_nxt_reg_10_11_inst : DLH_X1 port map( G => n27538, D => n27338, Q => 
                           regs_nxt_10_11_port);
   regs_reg_10_11_inst : DFF_X1 port map( D => N706, CK => clk, Q => n_1325, QN
                           => n25302);
   regs_nxt_reg_10_10_inst : DLH_X1 port map( G => n27538, D => n27344, Q => 
                           regs_nxt_10_10_port);
   regs_reg_10_10_inst : DFF_X1 port map( D => N705, CK => clk, Q => n_1326, QN
                           => n25301);
   regs_nxt_reg_10_9_inst : DLH_X1 port map( G => n27539, D => n27350, Q => 
                           regs_nxt_10_9_port);
   regs_reg_10_9_inst : DFF_X1 port map( D => N704, CK => clk, Q => n_1327, QN 
                           => n25300);
   regs_nxt_reg_10_8_inst : DLH_X1 port map( G => n27539, D => n27356, Q => 
                           regs_nxt_10_8_port);
   regs_reg_10_8_inst : DFF_X1 port map( D => N703, CK => clk, Q => n_1328, QN 
                           => n25299);
   regs_nxt_reg_10_7_inst : DLH_X1 port map( G => n27539, D => n27362, Q => 
                           regs_nxt_10_7_port);
   regs_reg_10_7_inst : DFF_X1 port map( D => N702, CK => clk, Q => n_1329, QN 
                           => n25298);
   regs_nxt_reg_10_6_inst : DLH_X1 port map( G => n27539, D => n27368, Q => 
                           regs_nxt_10_6_port);
   regs_reg_10_6_inst : DFF_X1 port map( D => N701, CK => clk, Q => n_1330, QN 
                           => n25297);
   regs_nxt_reg_10_5_inst : DLH_X1 port map( G => n27539, D => n27278, Q => 
                           regs_nxt_10_5_port);
   regs_reg_10_5_inst : DFF_X1 port map( D => N700, CK => clk, Q => n_1331, QN 
                           => n25296);
   regs_nxt_reg_10_4_inst : DLH_X1 port map( G => n27539, D => n27440, Q => 
                           regs_nxt_10_4_port);
   regs_reg_10_4_inst : DFF_X1 port map( D => N699, CK => clk, Q => n_1332, QN 
                           => n25295);
   regs_nxt_reg_10_3_inst : DLH_X1 port map( G => n27540, D => n27446, Q => 
                           regs_nxt_10_3_port);
   regs_reg_10_3_inst : DFF_X1 port map( D => N698, CK => clk, Q => n_1333, QN 
                           => n25294);
   regs_nxt_reg_10_2_inst : DLH_X1 port map( G => n27539, D => n27452, Q => 
                           regs_nxt_10_2_port);
   regs_reg_10_2_inst : DFF_X1 port map( D => N697, CK => clk, Q => n_1334, QN 
                           => n25293);
   regs_nxt_reg_10_1_inst : DLH_X1 port map( G => n27538, D => n27458, Q => 
                           regs_nxt_10_1_port);
   regs_reg_10_1_inst : DFF_X1 port map( D => N696, CK => clk, Q => n_1335, QN 
                           => n25292);
   regs_nxt_reg_10_0_inst : DLH_X1 port map( G => n27539, D => n27464, Q => 
                           regs_nxt_10_0_port);
   regs_reg_10_0_inst : DFF_X1 port map( D => N695, CK => clk, Q => n_1336, QN 
                           => n25291);
   regs_nxt_reg_11_31_inst : DLH_X1 port map( G => n27546, D => n27374, Q => 
                           regs_nxt_11_31_port);
   regs_reg_11_31_inst : DFF_X1 port map( D => N694, CK => clk, Q => n25244, QN
                           => n_1337);
   regs_nxt_reg_11_30_inst : DLH_X1 port map( G => n27546, D => n27380, Q => 
                           regs_nxt_11_30_port);
   regs_reg_11_30_inst : DFF_X1 port map( D => N693, CK => clk, Q => n25243, QN
                           => n_1338);
   regs_nxt_reg_11_29_inst : DLH_X1 port map( G => n27545, D => n27386, Q => 
                           regs_nxt_11_29_port);
   regs_reg_11_29_inst : DFF_X1 port map( D => N692, CK => clk, Q => n25242, QN
                           => n_1339);
   regs_nxt_reg_11_28_inst : DLH_X1 port map( G => n27545, D => n27392, Q => 
                           regs_nxt_11_28_port);
   regs_reg_11_28_inst : DFF_X1 port map( D => N691, CK => clk, Q => n25241, QN
                           => n_1340);
   regs_nxt_reg_11_27_inst : DLH_X1 port map( G => n27548, D => n27398, Q => 
                           regs_nxt_11_27_port);
   regs_reg_11_27_inst : DFF_X1 port map( D => N690, CK => clk, Q => n25240, QN
                           => n_1341);
   regs_nxt_reg_11_26_inst : DLH_X1 port map( G => n27547, D => n27404, Q => 
                           regs_nxt_11_26_port);
   regs_reg_11_26_inst : DFF_X1 port map( D => N689, CK => clk, Q => n25239, QN
                           => n_1342);
   regs_nxt_reg_11_25_inst : DLH_X1 port map( G => n27548, D => n27410, Q => 
                           regs_nxt_11_25_port);
   regs_reg_11_25_inst : DFF_X1 port map( D => N688, CK => clk, Q => n25238, QN
                           => n_1343);
   regs_nxt_reg_11_24_inst : DLH_X1 port map( G => n27547, D => n27416, Q => 
                           regs_nxt_11_24_port);
   regs_reg_11_24_inst : DFF_X1 port map( D => N687, CK => clk, Q => n25237, QN
                           => n_1344);
   regs_nxt_reg_11_23_inst : DLH_X1 port map( G => n27547, D => n27422, Q => 
                           regs_nxt_11_23_port);
   regs_reg_11_23_inst : DFF_X1 port map( D => N686, CK => clk, Q => n25236, QN
                           => n_1345);
   regs_nxt_reg_11_22_inst : DLH_X1 port map( G => n27547, D => n27428, Q => 
                           regs_nxt_11_22_port);
   regs_reg_11_22_inst : DFF_X1 port map( D => N685, CK => clk, Q => n26752, QN
                           => n2358);
   regs_nxt_reg_11_21_inst : DLH_X1 port map( G => n27545, D => n27434, Q => 
                           regs_nxt_11_21_port);
   regs_reg_11_21_inst : DFF_X1 port map( D => N684, CK => clk, Q => n26751, QN
                           => n2354);
   regs_nxt_reg_11_20_inst : DLH_X1 port map( G => n27545, D => n27284, Q => 
                           regs_nxt_11_20_port);
   regs_reg_11_20_inst : DFF_X1 port map( D => N683, CK => clk, Q => n26750, QN
                           => n2350);
   regs_nxt_reg_11_19_inst : DLH_X1 port map( G => n27545, D => n27290, Q => 
                           regs_nxt_11_19_port);
   regs_reg_11_19_inst : DFF_X1 port map( D => N682, CK => clk, Q => n26749, QN
                           => n2346);
   regs_nxt_reg_11_18_inst : DLH_X1 port map( G => n27547, D => n27296, Q => 
                           regs_nxt_11_18_port);
   regs_reg_11_18_inst : DFF_X1 port map( D => N681, CK => clk, Q => n26748, QN
                           => n2342);
   regs_nxt_reg_11_17_inst : DLH_X1 port map( G => n27545, D => n27302, Q => 
                           regs_nxt_11_17_port);
   regs_reg_11_17_inst : DFF_X1 port map( D => N680, CK => clk, Q => n26747, QN
                           => n2338);
   regs_nxt_reg_11_16_inst : DLH_X1 port map( G => n27547, D => n27308, Q => 
                           regs_nxt_11_16_port);
   regs_reg_11_16_inst : DFF_X1 port map( D => N679, CK => clk, Q => n26746, QN
                           => n2334);
   regs_nxt_reg_11_15_inst : DLH_X1 port map( G => n27545, D => n27314, Q => 
                           regs_nxt_11_15_port);
   regs_reg_11_15_inst : DFF_X1 port map( D => N678, CK => clk, Q => n26745, QN
                           => n2330);
   regs_nxt_reg_11_14_inst : DLH_X1 port map( G => n27547, D => n27320, Q => 
                           regs_nxt_11_14_port);
   regs_reg_11_14_inst : DFF_X1 port map( D => N677, CK => clk, Q => n26744, QN
                           => n2326);
   regs_nxt_reg_11_13_inst : DLH_X1 port map( G => n27547, D => n27326, Q => 
                           regs_nxt_11_13_port);
   regs_reg_11_13_inst : DFF_X1 port map( D => N676, CK => clk, Q => n26743, QN
                           => n2322);
   regs_nxt_reg_11_12_inst : DLH_X1 port map( G => n27547, D => n27332, Q => 
                           regs_nxt_11_12_port);
   regs_reg_11_12_inst : DFF_X1 port map( D => N675, CK => clk, Q => n26742, QN
                           => n2318);
   regs_nxt_reg_11_11_inst : DLH_X1 port map( G => n27545, D => n27338, Q => 
                           regs_nxt_11_11_port);
   regs_reg_11_11_inst : DFF_X1 port map( D => N674, CK => clk, Q => n26741, QN
                           => n2314);
   regs_nxt_reg_11_10_inst : DLH_X1 port map( G => n27545, D => n27344, Q => 
                           regs_nxt_11_10_port);
   regs_reg_11_10_inst : DFF_X1 port map( D => N673, CK => clk, Q => n26740, QN
                           => n2310);
   regs_nxt_reg_11_9_inst : DLH_X1 port map( G => n27546, D => n27350, Q => 
                           regs_nxt_11_9_port);
   regs_reg_11_9_inst : DFF_X1 port map( D => N672, CK => clk, Q => n26739, QN 
                           => n2306);
   regs_nxt_reg_11_8_inst : DLH_X1 port map( G => n27546, D => n27356, Q => 
                           regs_nxt_11_8_port);
   regs_reg_11_8_inst : DFF_X1 port map( D => N671, CK => clk, Q => n26738, QN 
                           => n2302);
   regs_nxt_reg_11_7_inst : DLH_X1 port map( G => n27546, D => n27362, Q => 
                           regs_nxt_11_7_port);
   regs_reg_11_7_inst : DFF_X1 port map( D => N670, CK => clk, Q => n26737, QN 
                           => n2298);
   regs_nxt_reg_11_6_inst : DLH_X1 port map( G => n27546, D => n27368, Q => 
                           regs_nxt_11_6_port);
   regs_reg_11_6_inst : DFF_X1 port map( D => N669, CK => clk, Q => n26736, QN 
                           => n2294);
   regs_nxt_reg_11_5_inst : DLH_X1 port map( G => n27546, D => n27278, Q => 
                           regs_nxt_11_5_port);
   regs_reg_11_5_inst : DFF_X1 port map( D => N668, CK => clk, Q => n26735, QN 
                           => n2290);
   regs_nxt_reg_11_4_inst : DLH_X1 port map( G => n27546, D => n27440, Q => 
                           regs_nxt_11_4_port);
   regs_reg_11_4_inst : DFF_X1 port map( D => N667, CK => clk, Q => n26734, QN 
                           => n2656);
   regs_nxt_reg_11_3_inst : DLH_X1 port map( G => n27547, D => n27446, Q => 
                           regs_nxt_11_3_port);
   regs_reg_11_3_inst : DFF_X1 port map( D => N666, CK => clk, Q => n26733, QN 
                           => n2654);
   regs_nxt_reg_11_2_inst : DLH_X1 port map( G => n27546, D => n27452, Q => 
                           regs_nxt_11_2_port);
   regs_reg_11_2_inst : DFF_X1 port map( D => N665, CK => clk, Q => n26732, QN 
                           => n2652);
   regs_nxt_reg_11_1_inst : DLH_X1 port map( G => n27545, D => n27458, Q => 
                           regs_nxt_11_1_port);
   regs_reg_11_1_inst : DFF_X1 port map( D => N664, CK => clk, Q => n26731, QN 
                           => n2650);
   regs_nxt_reg_11_0_inst : DLH_X1 port map( G => n27546, D => n27464, Q => 
                           regs_nxt_11_0_port);
   regs_reg_11_0_inst : DFF_X1 port map( D => N663, CK => clk, Q => n26730, QN 
                           => n2648);
   regs_nxt_reg_12_31_inst : DLH_X1 port map( G => n27553, D => n27374, Q => 
                           regs_nxt_12_31_port);
   regs_reg_12_31_inst : DFF_X1 port map( D => N662, CK => clk, Q => n_1346, QN
                           => n25258);
   regs_nxt_reg_12_30_inst : DLH_X1 port map( G => n27553, D => n27380, Q => 
                           regs_nxt_12_30_port);
   regs_reg_12_30_inst : DFF_X1 port map( D => N661, CK => clk, Q => n_1347, QN
                           => n25257);
   regs_nxt_reg_12_29_inst : DLH_X1 port map( G => n27554, D => n27386, Q => 
                           regs_nxt_12_29_port);
   regs_reg_12_29_inst : DFF_X1 port map( D => N660, CK => clk, Q => n_1348, QN
                           => n25256);
   regs_nxt_reg_12_28_inst : DLH_X1 port map( G => n27552, D => n27392, Q => 
                           regs_nxt_12_28_port);
   regs_reg_12_28_inst : DFF_X1 port map( D => N659, CK => clk, Q => n_1349, QN
                           => n25255);
   regs_nxt_reg_12_27_inst : DLH_X1 port map( G => n27555, D => n27398, Q => 
                           regs_nxt_12_27_port);
   regs_reg_12_27_inst : DFF_X1 port map( D => N658, CK => clk, Q => n_1350, QN
                           => n25254);
   regs_nxt_reg_12_26_inst : DLH_X1 port map( G => n27554, D => n27404, Q => 
                           regs_nxt_12_26_port);
   regs_reg_12_26_inst : DFF_X1 port map( D => N657, CK => clk, Q => n_1351, QN
                           => n25253);
   regs_nxt_reg_12_25_inst : DLH_X1 port map( G => n27555, D => n27410, Q => 
                           regs_nxt_12_25_port);
   regs_reg_12_25_inst : DFF_X1 port map( D => N656, CK => clk, Q => n_1352, QN
                           => n25252);
   regs_nxt_reg_12_24_inst : DLH_X1 port map( G => n27554, D => n27416, Q => 
                           regs_nxt_12_24_port);
   regs_reg_12_24_inst : DFF_X1 port map( D => N655, CK => clk, Q => n_1353, QN
                           => n25251);
   regs_nxt_reg_12_23_inst : DLH_X1 port map( G => n27552, D => n27422, Q => 
                           regs_nxt_12_23_port);
   regs_reg_12_23_inst : DFF_X1 port map( D => N654, CK => clk, Q => n_1354, QN
                           => n25250);
   regs_nxt_reg_12_22_inst : DLH_X1 port map( G => n27554, D => n27428, Q => 
                           regs_nxt_12_22_port);
   regs_reg_12_22_inst : DFF_X1 port map( D => N653, CK => clk, Q => n2356, QN 
                           => n26929);
   regs_nxt_reg_12_21_inst : DLH_X1 port map( G => n27552, D => n27434, Q => 
                           regs_nxt_12_21_port);
   regs_reg_12_21_inst : DFF_X1 port map( D => N652, CK => clk, Q => n2352, QN 
                           => n26928);
   regs_nxt_reg_12_20_inst : DLH_X1 port map( G => n27552, D => n27284, Q => 
                           regs_nxt_12_20_port);
   regs_reg_12_20_inst : DFF_X1 port map( D => N651, CK => clk, Q => n2348, QN 
                           => n26927);
   regs_nxt_reg_12_19_inst : DLH_X1 port map( G => n27552, D => n27290, Q => 
                           regs_nxt_12_19_port);
   regs_reg_12_19_inst : DFF_X1 port map( D => N650, CK => clk, Q => n2344, QN 
                           => n26926);
   regs_nxt_reg_12_18_inst : DLH_X1 port map( G => n27554, D => n27296, Q => 
                           regs_nxt_12_18_port);
   regs_reg_12_18_inst : DFF_X1 port map( D => N649, CK => clk, Q => n2340, QN 
                           => n26925);
   regs_nxt_reg_12_17_inst : DLH_X1 port map( G => n27552, D => n27302, Q => 
                           regs_nxt_12_17_port);
   regs_reg_12_17_inst : DFF_X1 port map( D => N648, CK => clk, Q => n2336, QN 
                           => n26924);
   regs_nxt_reg_12_16_inst : DLH_X1 port map( G => n27554, D => n27308, Q => 
                           regs_nxt_12_16_port);
   regs_reg_12_16_inst : DFF_X1 port map( D => N647, CK => clk, Q => n2332, QN 
                           => n26923);
   regs_nxt_reg_12_15_inst : DLH_X1 port map( G => n27552, D => n27314, Q => 
                           regs_nxt_12_15_port);
   regs_reg_12_15_inst : DFF_X1 port map( D => N646, CK => clk, Q => n2328, QN 
                           => n26922);
   regs_nxt_reg_12_14_inst : DLH_X1 port map( G => n27554, D => n27320, Q => 
                           regs_nxt_12_14_port);
   regs_reg_12_14_inst : DFF_X1 port map( D => N645, CK => clk, Q => n2324, QN 
                           => n26921);
   regs_nxt_reg_12_13_inst : DLH_X1 port map( G => n27552, D => n27326, Q => 
                           regs_nxt_12_13_port);
   regs_reg_12_13_inst : DFF_X1 port map( D => N644, CK => clk, Q => n2320, QN 
                           => n26920);
   regs_nxt_reg_12_12_inst : DLH_X1 port map( G => n27554, D => n27332, Q => 
                           regs_nxt_12_12_port);
   regs_reg_12_12_inst : DFF_X1 port map( D => N643, CK => clk, Q => n2316, QN 
                           => n26919);
   regs_nxt_reg_12_11_inst : DLH_X1 port map( G => n27552, D => n27338, Q => 
                           regs_nxt_12_11_port);
   regs_reg_12_11_inst : DFF_X1 port map( D => N642, CK => clk, Q => n2312, QN 
                           => n26918);
   regs_nxt_reg_12_10_inst : DLH_X1 port map( G => n27554, D => n27344, Q => 
                           regs_nxt_12_10_port);
   regs_reg_12_10_inst : DFF_X1 port map( D => N641, CK => clk, Q => n2308, QN 
                           => n26917);
   regs_nxt_reg_12_9_inst : DLH_X1 port map( G => n27553, D => n27350, Q => 
                           regs_nxt_12_9_port);
   regs_reg_12_9_inst : DFF_X1 port map( D => N640, CK => clk, Q => n2304, QN 
                           => n26916);
   regs_nxt_reg_12_8_inst : DLH_X1 port map( G => n27553, D => n27356, Q => 
                           regs_nxt_12_8_port);
   regs_reg_12_8_inst : DFF_X1 port map( D => N639, CK => clk, Q => n2300, QN 
                           => n26915);
   regs_nxt_reg_12_7_inst : DLH_X1 port map( G => n27553, D => n27362, Q => 
                           regs_nxt_12_7_port);
   regs_reg_12_7_inst : DFF_X1 port map( D => N638, CK => clk, Q => n2296, QN 
                           => n26914);
   regs_nxt_reg_12_6_inst : DLH_X1 port map( G => n27553, D => n27368, Q => 
                           regs_nxt_12_6_port);
   regs_reg_12_6_inst : DFF_X1 port map( D => N637, CK => clk, Q => n2292, QN 
                           => n26913);
   regs_nxt_reg_12_5_inst : DLH_X1 port map( G => n27553, D => n27278, Q => 
                           regs_nxt_12_5_port);
   regs_reg_12_5_inst : DFF_X1 port map( D => N636, CK => clk, Q => n2288, QN 
                           => n26912);
   regs_nxt_reg_12_4_inst : DLH_X1 port map( G => n27553, D => n27440, Q => 
                           regs_nxt_12_4_port);
   regs_reg_12_4_inst : DFF_X1 port map( D => N635, CK => clk, Q => n2647_port,
                           QN => n26911);
   regs_nxt_reg_12_3_inst : DLH_X1 port map( G => n27554, D => n27444, Q => 
                           regs_nxt_12_3_port);
   regs_reg_12_3_inst : DFF_X1 port map( D => N634, CK => clk, Q => n2645, QN 
                           => n26910);
   regs_nxt_reg_12_2_inst : DLH_X1 port map( G => n27553, D => n27450, Q => 
                           regs_nxt_12_2_port);
   regs_reg_12_2_inst : DFF_X1 port map( D => N633, CK => clk, Q => n2643, QN 
                           => n26909);
   regs_nxt_reg_12_1_inst : DLH_X1 port map( G => n27552, D => n27458, Q => 
                           regs_nxt_12_1_port);
   regs_reg_12_1_inst : DFF_X1 port map( D => N632, CK => clk, Q => n2641, QN 
                           => n26908);
   regs_nxt_reg_12_0_inst : DLH_X1 port map( G => n27553, D => n27464, Q => 
                           regs_nxt_12_0_port);
   regs_reg_12_0_inst : DFF_X1 port map( D => N631, CK => clk, Q => n2639, QN 
                           => n26907);
   regs_nxt_reg_13_31_inst : DLH_X1 port map( G => n27560, D => n27374, Q => 
                           regs_nxt_13_31_port);
   regs_reg_13_31_inst : DFF_X1 port map( D => N630, CK => clk, Q => 
                           regs_13_31_port, QN => n_1355);
   regs_nxt_reg_13_30_inst : DLH_X1 port map( G => n27560, D => n27380, Q => 
                           regs_nxt_13_30_port);
   regs_reg_13_30_inst : DFF_X1 port map( D => N629, CK => clk, Q => 
                           regs_13_30_port, QN => n_1356);
   regs_nxt_reg_13_29_inst : DLH_X1 port map( G => n27559, D => n27386, Q => 
                           regs_nxt_13_29_port);
   regs_reg_13_29_inst : DFF_X1 port map( D => N628, CK => clk, Q => 
                           regs_13_29_port, QN => n_1357);
   regs_nxt_reg_13_28_inst : DLH_X1 port map( G => n27559, D => n27392, Q => 
                           regs_nxt_13_28_port);
   regs_reg_13_28_inst : DFF_X1 port map( D => N627, CK => clk, Q => 
                           regs_13_28_port, QN => n_1358);
   regs_nxt_reg_13_27_inst : DLH_X1 port map( G => n27562, D => n27398, Q => 
                           regs_nxt_13_27_port);
   regs_reg_13_27_inst : DFF_X1 port map( D => N626, CK => clk, Q => 
                           regs_13_27_port, QN => n_1359);
   regs_nxt_reg_13_26_inst : DLH_X1 port map( G => n27561, D => n27404, Q => 
                           regs_nxt_13_26_port);
   regs_reg_13_26_inst : DFF_X1 port map( D => N625, CK => clk, Q => 
                           regs_13_26_port, QN => n_1360);
   regs_nxt_reg_13_25_inst : DLH_X1 port map( G => n27562, D => n27410, Q => 
                           regs_nxt_13_25_port);
   regs_reg_13_25_inst : DFF_X1 port map( D => N624, CK => clk, Q => 
                           regs_13_25_port, QN => n_1361);
   regs_nxt_reg_13_24_inst : DLH_X1 port map( G => n27561, D => n27416, Q => 
                           regs_nxt_13_24_port);
   regs_reg_13_24_inst : DFF_X1 port map( D => N623, CK => clk, Q => 
                           regs_13_24_port, QN => n_1362);
   regs_nxt_reg_13_23_inst : DLH_X1 port map( G => n27561, D => n27422, Q => 
                           regs_nxt_13_23_port);
   regs_reg_13_23_inst : DFF_X1 port map( D => N622, CK => clk, Q => 
                           regs_13_23_port, QN => n_1363);
   regs_nxt_reg_13_22_inst : DLH_X1 port map( G => n27561, D => n27428, Q => 
                           regs_nxt_13_22_port);
   regs_reg_13_22_inst : DFF_X1 port map( D => N621, CK => clk, Q => 
                           regs_13_22_port, QN => n_1364);
   regs_nxt_reg_13_21_inst : DLH_X1 port map( G => n27559, D => n27434, Q => 
                           regs_nxt_13_21_port);
   regs_reg_13_21_inst : DFF_X1 port map( D => N620, CK => clk, Q => 
                           regs_13_21_port, QN => n_1365);
   regs_nxt_reg_13_20_inst : DLH_X1 port map( G => n27559, D => n27284, Q => 
                           regs_nxt_13_20_port);
   regs_reg_13_20_inst : DFF_X1 port map( D => N619, CK => clk, Q => 
                           regs_13_20_port, QN => n_1366);
   regs_nxt_reg_13_19_inst : DLH_X1 port map( G => n27559, D => n27290, Q => 
                           regs_nxt_13_19_port);
   regs_reg_13_19_inst : DFF_X1 port map( D => N618, CK => clk, Q => 
                           regs_13_19_port, QN => n_1367);
   regs_nxt_reg_13_18_inst : DLH_X1 port map( G => n27561, D => n27296, Q => 
                           regs_nxt_13_18_port);
   regs_reg_13_18_inst : DFF_X1 port map( D => N617, CK => clk, Q => 
                           regs_13_18_port, QN => n_1368);
   regs_nxt_reg_13_17_inst : DLH_X1 port map( G => n27559, D => n27302, Q => 
                           regs_nxt_13_17_port);
   regs_reg_13_17_inst : DFF_X1 port map( D => N616, CK => clk, Q => 
                           regs_13_17_port, QN => n_1369);
   regs_nxt_reg_13_16_inst : DLH_X1 port map( G => n27561, D => n27308, Q => 
                           regs_nxt_13_16_port);
   regs_reg_13_16_inst : DFF_X1 port map( D => N615, CK => clk, Q => 
                           regs_13_16_port, QN => n_1370);
   regs_nxt_reg_13_15_inst : DLH_X1 port map( G => n27559, D => n27314, Q => 
                           regs_nxt_13_15_port);
   regs_reg_13_15_inst : DFF_X1 port map( D => N614, CK => clk, Q => 
                           regs_13_15_port, QN => n_1371);
   regs_nxt_reg_13_14_inst : DLH_X1 port map( G => n27561, D => n27320, Q => 
                           regs_nxt_13_14_port);
   regs_reg_13_14_inst : DFF_X1 port map( D => N613, CK => clk, Q => 
                           regs_13_14_port, QN => n_1372);
   regs_nxt_reg_13_13_inst : DLH_X1 port map( G => n27561, D => n27326, Q => 
                           regs_nxt_13_13_port);
   regs_reg_13_13_inst : DFF_X1 port map( D => N612, CK => clk, Q => 
                           regs_13_13_port, QN => n_1373);
   regs_nxt_reg_13_12_inst : DLH_X1 port map( G => n27561, D => n27332, Q => 
                           regs_nxt_13_12_port);
   regs_reg_13_12_inst : DFF_X1 port map( D => N611, CK => clk, Q => 
                           regs_13_12_port, QN => n_1374);
   regs_nxt_reg_13_11_inst : DLH_X1 port map( G => n27559, D => n27338, Q => 
                           regs_nxt_13_11_port);
   regs_reg_13_11_inst : DFF_X1 port map( D => N610, CK => clk, Q => 
                           regs_13_11_port, QN => n_1375);
   regs_nxt_reg_13_10_inst : DLH_X1 port map( G => n27559, D => n27344, Q => 
                           regs_nxt_13_10_port);
   regs_reg_13_10_inst : DFF_X1 port map( D => N609, CK => clk, Q => 
                           regs_13_10_port, QN => n_1376);
   regs_nxt_reg_13_9_inst : DLH_X1 port map( G => n27560, D => n27350, Q => 
                           regs_nxt_13_9_port);
   regs_reg_13_9_inst : DFF_X1 port map( D => N608, CK => clk, Q => 
                           regs_13_9_port, QN => n_1377);
   regs_nxt_reg_13_8_inst : DLH_X1 port map( G => n27560, D => n27356, Q => 
                           regs_nxt_13_8_port);
   regs_reg_13_8_inst : DFF_X1 port map( D => N607, CK => clk, Q => 
                           regs_13_8_port, QN => n_1378);
   regs_nxt_reg_13_7_inst : DLH_X1 port map( G => n27560, D => n27362, Q => 
                           regs_nxt_13_7_port);
   regs_reg_13_7_inst : DFF_X1 port map( D => N606, CK => clk, Q => 
                           regs_13_7_port, QN => n_1379);
   regs_nxt_reg_13_6_inst : DLH_X1 port map( G => n27560, D => n27368, Q => 
                           regs_nxt_13_6_port);
   regs_reg_13_6_inst : DFF_X1 port map( D => N605, CK => clk, Q => 
                           regs_13_6_port, QN => n_1380);
   regs_nxt_reg_13_5_inst : DLH_X1 port map( G => n27560, D => n27278, Q => 
                           regs_nxt_13_5_port);
   regs_reg_13_5_inst : DFF_X1 port map( D => N604, CK => clk, Q => 
                           regs_13_5_port, QN => n_1381);
   regs_nxt_reg_13_4_inst : DLH_X1 port map( G => n27560, D => n27440, Q => 
                           regs_nxt_13_4_port);
   regs_reg_13_4_inst : DFF_X1 port map( D => N603, CK => clk, Q => 
                           regs_13_4_port, QN => n_1382);
   regs_nxt_reg_13_3_inst : DLH_X1 port map( G => n27561, D => n27446, Q => 
                           regs_nxt_13_3_port);
   regs_reg_13_3_inst : DFF_X1 port map( D => N602, CK => clk, Q => 
                           regs_13_3_port, QN => n_1383);
   regs_nxt_reg_13_2_inst : DLH_X1 port map( G => n27560, D => n27452, Q => 
                           regs_nxt_13_2_port);
   regs_reg_13_2_inst : DFF_X1 port map( D => N601, CK => clk, Q => 
                           regs_13_2_port, QN => n_1384);
   regs_nxt_reg_13_1_inst : DLH_X1 port map( G => n27559, D => n27458, Q => 
                           regs_nxt_13_1_port);
   regs_reg_13_1_inst : DFF_X1 port map( D => N600, CK => clk, Q => 
                           regs_13_1_port, QN => n_1385);
   regs_nxt_reg_13_0_inst : DLH_X1 port map( G => n27560, D => n27464, Q => 
                           regs_nxt_13_0_port);
   regs_reg_13_0_inst : DFF_X1 port map( D => N599, CK => clk, Q => 
                           regs_13_0_port, QN => n_1386);
   regs_nxt_reg_14_31_inst : DLH_X1 port map( G => n27567, D => n27374, Q => 
                           regs_nxt_14_31_port);
   regs_reg_14_31_inst : DFF_X1 port map( D => N598, CK => clk, Q => n26764, QN
                           => n2219);
   regs_nxt_reg_14_30_inst : DLH_X1 port map( G => n27567, D => n27380, Q => 
                           regs_nxt_14_30_port);
   regs_reg_14_30_inst : DFF_X1 port map( D => N597, CK => clk, Q => n26763, QN
                           => n2212);
   regs_nxt_reg_14_29_inst : DLH_X1 port map( G => n27568, D => n27386, Q => 
                           regs_nxt_14_29_port);
   regs_reg_14_29_inst : DFF_X1 port map( D => N596, CK => clk, Q => n26762, QN
                           => n2205);
   regs_nxt_reg_14_28_inst : DLH_X1 port map( G => n27566, D => n27392, Q => 
                           regs_nxt_14_28_port);
   regs_reg_14_28_inst : DFF_X1 port map( D => N595, CK => clk, Q => n26761, QN
                           => n2198);
   regs_nxt_reg_14_27_inst : DLH_X1 port map( G => n27568, D => n27398, Q => 
                           regs_nxt_14_27_port);
   regs_reg_14_27_inst : DFF_X1 port map( D => N594, CK => clk, Q => n26760, QN
                           => n2191);
   regs_nxt_reg_14_26_inst : DLH_X1 port map( G => n27568, D => n27404, Q => 
                           regs_nxt_14_26_port);
   regs_reg_14_26_inst : DFF_X1 port map( D => N593, CK => clk, Q => n26759, QN
                           => n2184);
   regs_nxt_reg_14_25_inst : DLH_X1 port map( G => n27569, D => n27410, Q => 
                           regs_nxt_14_25_port);
   regs_reg_14_25_inst : DFF_X1 port map( D => N592, CK => clk, Q => n26758, QN
                           => n2177);
   regs_nxt_reg_14_24_inst : DLH_X1 port map( G => n27568, D => n27416, Q => 
                           regs_nxt_14_24_port);
   regs_reg_14_24_inst : DFF_X1 port map( D => N591, CK => clk, Q => n26757, QN
                           => n2170);
   regs_nxt_reg_14_23_inst : DLH_X1 port map( G => n27569, D => n27422, Q => 
                           regs_nxt_14_23_port);
   regs_reg_14_23_inst : DFF_X1 port map( D => N590, CK => clk, Q => n26756, QN
                           => n2163);
   regs_nxt_reg_14_22_inst : DLH_X1 port map( G => n27568, D => n27428, Q => 
                           regs_nxt_14_22_port);
   regs_reg_14_22_inst : DFF_X1 port map( D => N589, CK => clk, Q => n26755, QN
                           => n2156);
   regs_nxt_reg_14_21_inst : DLH_X1 port map( G => n27566, D => n27434, Q => 
                           regs_nxt_14_21_port);
   regs_reg_14_21_inst : DFF_X1 port map( D => N588, CK => clk, Q => n26754, QN
                           => n2149);
   regs_nxt_reg_14_20_inst : DLH_X1 port map( G => n27566, D => n27284, Q => 
                           regs_nxt_14_20_port);
   regs_reg_14_20_inst : DFF_X1 port map( D => N587, CK => clk, Q => n26753, QN
                           => n2142);
   regs_nxt_reg_14_19_inst : DLH_X1 port map( G => n27566, D => n27290, Q => 
                           regs_nxt_14_19_port);
   regs_reg_14_19_inst : DFF_X1 port map( D => N586, CK => clk, Q => n25230, QN
                           => n_1387);
   regs_nxt_reg_14_18_inst : DLH_X1 port map( G => n27568, D => n27296, Q => 
                           regs_nxt_14_18_port);
   regs_reg_14_18_inst : DFF_X1 port map( D => N585, CK => clk, Q => n25229, QN
                           => n_1388);
   regs_nxt_reg_14_17_inst : DLH_X1 port map( G => n27566, D => n27302, Q => 
                           regs_nxt_14_17_port);
   regs_reg_14_17_inst : DFF_X1 port map( D => N584, CK => clk, Q => n25228, QN
                           => n_1389);
   regs_nxt_reg_14_16_inst : DLH_X1 port map( G => n27568, D => n27308, Q => 
                           regs_nxt_14_16_port);
   regs_reg_14_16_inst : DFF_X1 port map( D => N583, CK => clk, Q => n25227, QN
                           => n_1390);
   regs_nxt_reg_14_15_inst : DLH_X1 port map( G => n27566, D => n27314, Q => 
                           regs_nxt_14_15_port);
   regs_reg_14_15_inst : DFF_X1 port map( D => N582, CK => clk, Q => n25226, QN
                           => n_1391);
   regs_nxt_reg_14_14_inst : DLH_X1 port map( G => n27568, D => n27320, Q => 
                           regs_nxt_14_14_port);
   regs_reg_14_14_inst : DFF_X1 port map( D => N581, CK => clk, Q => n25225, QN
                           => n_1392);
   regs_nxt_reg_14_13_inst : DLH_X1 port map( G => n27566, D => n27326, Q => 
                           regs_nxt_14_13_port);
   regs_reg_14_13_inst : DFF_X1 port map( D => N580, CK => clk, Q => n25224, QN
                           => n_1393);
   regs_nxt_reg_14_12_inst : DLH_X1 port map( G => n27568, D => n27332, Q => 
                           regs_nxt_14_12_port);
   regs_reg_14_12_inst : DFF_X1 port map( D => N579, CK => clk, Q => n25223, QN
                           => n_1394);
   regs_nxt_reg_14_11_inst : DLH_X1 port map( G => n27566, D => n27338, Q => 
                           regs_nxt_14_11_port);
   regs_reg_14_11_inst : DFF_X1 port map( D => N578, CK => clk, Q => n25222, QN
                           => n_1395);
   regs_nxt_reg_14_10_inst : DLH_X1 port map( G => n27566, D => n27344, Q => 
                           regs_nxt_14_10_port);
   regs_reg_14_10_inst : DFF_X1 port map( D => N577, CK => clk, Q => n25221, QN
                           => n_1396);
   regs_nxt_reg_14_9_inst : DLH_X1 port map( G => n27567, D => n27350, Q => 
                           regs_nxt_14_9_port);
   regs_reg_14_9_inst : DFF_X1 port map( D => N576, CK => clk, Q => n25220, QN 
                           => n_1397);
   regs_nxt_reg_14_8_inst : DLH_X1 port map( G => n27567, D => n27356, Q => 
                           regs_nxt_14_8_port);
   regs_reg_14_8_inst : DFF_X1 port map( D => N575, CK => clk, Q => n25219, QN 
                           => n_1398);
   regs_nxt_reg_14_7_inst : DLH_X1 port map( G => n27567, D => n27362, Q => 
                           regs_nxt_14_7_port);
   regs_reg_14_7_inst : DFF_X1 port map( D => N574, CK => clk, Q => n25218, QN 
                           => n_1399);
   regs_nxt_reg_14_6_inst : DLH_X1 port map( G => n27567, D => n27368, Q => 
                           regs_nxt_14_6_port);
   regs_reg_14_6_inst : DFF_X1 port map( D => N573, CK => clk, Q => n25217, QN 
                           => n_1400);
   regs_nxt_reg_14_5_inst : DLH_X1 port map( G => n27567, D => n27278, Q => 
                           regs_nxt_14_5_port);
   regs_reg_14_5_inst : DFF_X1 port map( D => N572, CK => clk, Q => n25216, QN 
                           => n_1401);
   regs_nxt_reg_14_4_inst : DLH_X1 port map( G => n27567, D => n27440, Q => 
                           regs_nxt_14_4_port);
   regs_reg_14_4_inst : DFF_X1 port map( D => N571, CK => clk, Q => n25215, QN 
                           => n_1402);
   regs_nxt_reg_14_3_inst : DLH_X1 port map( G => n27568, D => n27444, Q => 
                           regs_nxt_14_3_port);
   regs_reg_14_3_inst : DFF_X1 port map( D => N570, CK => clk, Q => n25214, QN 
                           => n_1403);
   regs_nxt_reg_14_2_inst : DLH_X1 port map( G => n27567, D => n27450, Q => 
                           regs_nxt_14_2_port);
   regs_reg_14_2_inst : DFF_X1 port map( D => N569, CK => clk, Q => n25213, QN 
                           => n_1404);
   regs_nxt_reg_14_1_inst : DLH_X1 port map( G => n27566, D => n27458, Q => 
                           regs_nxt_14_1_port);
   regs_reg_14_1_inst : DFF_X1 port map( D => N568, CK => clk, Q => n25212, QN 
                           => n_1405);
   regs_nxt_reg_14_0_inst : DLH_X1 port map( G => n27567, D => n27464, Q => 
                           regs_nxt_14_0_port);
   regs_reg_14_0_inst : DFF_X1 port map( D => N567, CK => clk, Q => n25211, QN 
                           => n_1406);
   regs_nxt_reg_15_31_inst : DLH_X1 port map( G => n27574, D => n27372, Q => 
                           regs_nxt_15_31_port);
   regs_reg_15_31_inst : DFF_X1 port map( D => N566, CK => clk, Q => 
                           regs_15_31_port, QN => n_1407);
   regs_nxt_reg_15_30_inst : DLH_X1 port map( G => n27574, D => n27378, Q => 
                           regs_nxt_15_30_port);
   regs_reg_15_30_inst : DFF_X1 port map( D => N565, CK => clk, Q => 
                           regs_15_30_port, QN => n_1408);
   regs_nxt_reg_15_29_inst : DLH_X1 port map( G => n27573, D => n27384, Q => 
                           regs_nxt_15_29_port);
   regs_reg_15_29_inst : DFF_X1 port map( D => N564, CK => clk, Q => 
                           regs_15_29_port, QN => n_1409);
   regs_nxt_reg_15_28_inst : DLH_X1 port map( G => n27573, D => n27390, Q => 
                           regs_nxt_15_28_port);
   regs_reg_15_28_inst : DFF_X1 port map( D => N563, CK => clk, Q => 
                           regs_15_28_port, QN => n_1410);
   regs_nxt_reg_15_27_inst : DLH_X1 port map( G => n27576, D => n27396, Q => 
                           regs_nxt_15_27_port);
   regs_reg_15_27_inst : DFF_X1 port map( D => N562, CK => clk, Q => 
                           regs_15_27_port, QN => n_1411);
   regs_nxt_reg_15_26_inst : DLH_X1 port map( G => n27575, D => n27402, Q => 
                           regs_nxt_15_26_port);
   regs_reg_15_26_inst : DFF_X1 port map( D => N561, CK => clk, Q => 
                           regs_15_26_port, QN => n_1412);
   regs_nxt_reg_15_25_inst : DLH_X1 port map( G => n27576, D => n27408, Q => 
                           regs_nxt_15_25_port);
   regs_reg_15_25_inst : DFF_X1 port map( D => N560, CK => clk, Q => 
                           regs_15_25_port, QN => n_1413);
   regs_nxt_reg_15_24_inst : DLH_X1 port map( G => n27575, D => n27414, Q => 
                           regs_nxt_15_24_port);
   regs_reg_15_24_inst : DFF_X1 port map( D => N559, CK => clk, Q => 
                           regs_15_24_port, QN => n_1414);
   regs_nxt_reg_15_23_inst : DLH_X1 port map( G => n27575, D => n27420, Q => 
                           regs_nxt_15_23_port);
   regs_reg_15_23_inst : DFF_X1 port map( D => N558, CK => clk, Q => 
                           regs_15_23_port, QN => n_1415);
   regs_nxt_reg_15_22_inst : DLH_X1 port map( G => n27575, D => n27426, Q => 
                           regs_nxt_15_22_port);
   regs_reg_15_22_inst : DFF_X1 port map( D => N557, CK => clk, Q => 
                           regs_15_22_port, QN => n_1416);
   regs_nxt_reg_15_21_inst : DLH_X1 port map( G => n27573, D => n27432, Q => 
                           regs_nxt_15_21_port);
   regs_reg_15_21_inst : DFF_X1 port map( D => N556, CK => clk, Q => 
                           regs_15_21_port, QN => n_1417);
   regs_nxt_reg_15_20_inst : DLH_X1 port map( G => n27573, D => n27282, Q => 
                           regs_nxt_15_20_port);
   regs_reg_15_20_inst : DFF_X1 port map( D => N555, CK => clk, Q => 
                           regs_15_20_port, QN => n_1418);
   regs_nxt_reg_15_19_inst : DLH_X1 port map( G => n27573, D => n27288, Q => 
                           regs_nxt_15_19_port);
   regs_reg_15_19_inst : DFF_X1 port map( D => N554, CK => clk, Q => 
                           regs_15_19_port, QN => n_1419);
   regs_nxt_reg_15_18_inst : DLH_X1 port map( G => n27575, D => n27294, Q => 
                           regs_nxt_15_18_port);
   regs_reg_15_18_inst : DFF_X1 port map( D => N553, CK => clk, Q => 
                           regs_15_18_port, QN => n_1420);
   regs_nxt_reg_15_17_inst : DLH_X1 port map( G => n27573, D => n27300, Q => 
                           regs_nxt_15_17_port);
   regs_reg_15_17_inst : DFF_X1 port map( D => N552, CK => clk, Q => 
                           regs_15_17_port, QN => n_1421);
   regs_nxt_reg_15_16_inst : DLH_X1 port map( G => n27575, D => n27306, Q => 
                           regs_nxt_15_16_port);
   regs_reg_15_16_inst : DFF_X1 port map( D => N551, CK => clk, Q => 
                           regs_15_16_port, QN => n_1422);
   regs_nxt_reg_15_15_inst : DLH_X1 port map( G => n27573, D => n27312, Q => 
                           regs_nxt_15_15_port);
   regs_reg_15_15_inst : DFF_X1 port map( D => N550, CK => clk, Q => 
                           regs_15_15_port, QN => n_1423);
   regs_nxt_reg_15_14_inst : DLH_X1 port map( G => n27575, D => n27318, Q => 
                           regs_nxt_15_14_port);
   regs_reg_15_14_inst : DFF_X1 port map( D => N549, CK => clk, Q => 
                           regs_15_14_port, QN => n_1424);
   regs_nxt_reg_15_13_inst : DLH_X1 port map( G => n27575, D => n27324, Q => 
                           regs_nxt_15_13_port);
   regs_reg_15_13_inst : DFF_X1 port map( D => N548, CK => clk, Q => 
                           regs_15_13_port, QN => n_1425);
   regs_nxt_reg_15_12_inst : DLH_X1 port map( G => n27575, D => n27330, Q => 
                           regs_nxt_15_12_port);
   regs_reg_15_12_inst : DFF_X1 port map( D => N547, CK => clk, Q => 
                           regs_15_12_port, QN => n_1426);
   regs_nxt_reg_15_11_inst : DLH_X1 port map( G => n27573, D => n27336, Q => 
                           regs_nxt_15_11_port);
   regs_reg_15_11_inst : DFF_X1 port map( D => N546, CK => clk, Q => 
                           regs_15_11_port, QN => n_1427);
   regs_nxt_reg_15_10_inst : DLH_X1 port map( G => n27573, D => n27342, Q => 
                           regs_nxt_15_10_port);
   regs_reg_15_10_inst : DFF_X1 port map( D => N545, CK => clk, Q => 
                           regs_15_10_port, QN => n_1428);
   regs_nxt_reg_15_9_inst : DLH_X1 port map( G => n27574, D => n27348, Q => 
                           regs_nxt_15_9_port);
   regs_reg_15_9_inst : DFF_X1 port map( D => N544, CK => clk, Q => 
                           regs_15_9_port, QN => n_1429);
   regs_nxt_reg_15_8_inst : DLH_X1 port map( G => n27574, D => n27354, Q => 
                           regs_nxt_15_8_port);
   regs_reg_15_8_inst : DFF_X1 port map( D => N543, CK => clk, Q => 
                           regs_15_8_port, QN => n_1430);
   regs_nxt_reg_15_7_inst : DLH_X1 port map( G => n27574, D => n27360, Q => 
                           regs_nxt_15_7_port);
   regs_reg_15_7_inst : DFF_X1 port map( D => N542, CK => clk, Q => 
                           regs_15_7_port, QN => n_1431);
   regs_nxt_reg_15_6_inst : DLH_X1 port map( G => n27574, D => n27366, Q => 
                           regs_nxt_15_6_port);
   regs_reg_15_6_inst : DFF_X1 port map( D => N541, CK => clk, Q => 
                           regs_15_6_port, QN => n_1432);
   regs_nxt_reg_15_5_inst : DLH_X1 port map( G => n27574, D => n27276, Q => 
                           regs_nxt_15_5_port);
   regs_reg_15_5_inst : DFF_X1 port map( D => N540, CK => clk, Q => 
                           regs_15_5_port, QN => n_1433);
   regs_nxt_reg_15_4_inst : DLH_X1 port map( G => n27574, D => n27438, Q => 
                           regs_nxt_15_4_port);
   regs_reg_15_4_inst : DFF_X1 port map( D => N539, CK => clk, Q => 
                           regs_15_4_port, QN => n_1434);
   regs_nxt_reg_15_3_inst : DLH_X1 port map( G => n27575, D => n27444, Q => 
                           regs_nxt_15_3_port);
   regs_reg_15_3_inst : DFF_X1 port map( D => N538, CK => clk, Q => 
                           regs_15_3_port, QN => n_1435);
   regs_nxt_reg_15_2_inst : DLH_X1 port map( G => n27574, D => n27450, Q => 
                           regs_nxt_15_2_port);
   regs_reg_15_2_inst : DFF_X1 port map( D => N537, CK => clk, Q => 
                           regs_15_2_port, QN => n_1436);
   regs_nxt_reg_15_1_inst : DLH_X1 port map( G => n27573, D => n27456, Q => 
                           regs_nxt_15_1_port);
   regs_reg_15_1_inst : DFF_X1 port map( D => N536, CK => clk, Q => 
                           regs_15_1_port, QN => n_1437);
   regs_nxt_reg_15_0_inst : DLH_X1 port map( G => n27574, D => n27462, Q => 
                           regs_nxt_15_0_port);
   regs_reg_15_0_inst : DFF_X1 port map( D => N535, CK => clk, Q => 
                           regs_15_0_port, QN => n_1438);
   regs_nxt_reg_16_31_inst : DLH_X1 port map( G => n27581, D => n27372, Q => 
                           regs_nxt_16_31_port);
   regs_reg_16_31_inst : DFF_X1 port map( D => N534, CK => clk, Q => n2012, QN 
                           => n26845);
   regs_nxt_reg_16_30_inst : DLH_X1 port map( G => n27581, D => n27378, Q => 
                           regs_nxt_16_30_port);
   regs_reg_16_30_inst : DFF_X1 port map( D => N533, CK => clk, Q => n2008, QN 
                           => n26844);
   regs_nxt_reg_16_29_inst : DLH_X1 port map( G => n27580, D => n27384, Q => 
                           regs_nxt_16_29_port);
   regs_reg_16_29_inst : DFF_X1 port map( D => N532, CK => clk, Q => n2004, QN 
                           => n26843);
   regs_nxt_reg_16_28_inst : DLH_X1 port map( G => n27580, D => n27390, Q => 
                           regs_nxt_16_28_port);
   regs_reg_16_28_inst : DFF_X1 port map( D => N531, CK => clk, Q => n2000, QN 
                           => n26842);
   regs_nxt_reg_16_27_inst : DLH_X1 port map( G => n27583, D => n27396, Q => 
                           regs_nxt_16_27_port);
   regs_reg_16_27_inst : DFF_X1 port map( D => N530, CK => clk, Q => n1996, QN 
                           => n26841);
   regs_nxt_reg_16_26_inst : DLH_X1 port map( G => n27582, D => n27402, Q => 
                           regs_nxt_16_26_port);
   regs_reg_16_26_inst : DFF_X1 port map( D => N529, CK => clk, Q => n1992, QN 
                           => n26840);
   regs_nxt_reg_16_25_inst : DLH_X1 port map( G => n27583, D => n27408, Q => 
                           regs_nxt_16_25_port);
   regs_reg_16_25_inst : DFF_X1 port map( D => N528, CK => clk, Q => n1988, QN 
                           => n26839);
   regs_nxt_reg_16_24_inst : DLH_X1 port map( G => n27582, D => n27414, Q => 
                           regs_nxt_16_24_port);
   regs_reg_16_24_inst : DFF_X1 port map( D => N527, CK => clk, Q => n1984, QN 
                           => n26838);
   regs_nxt_reg_16_23_inst : DLH_X1 port map( G => n27582, D => n27420, Q => 
                           regs_nxt_16_23_port);
   regs_reg_16_23_inst : DFF_X1 port map( D => N526, CK => clk, Q => n1980, QN 
                           => n26837);
   regs_nxt_reg_16_22_inst : DLH_X1 port map( G => n27582, D => n27426, Q => 
                           regs_nxt_16_22_port);
   regs_reg_16_22_inst : DFF_X1 port map( D => N525, CK => clk, Q => n1976, QN 
                           => n26836);
   regs_nxt_reg_16_21_inst : DLH_X1 port map( G => n27580, D => n27432, Q => 
                           regs_nxt_16_21_port);
   regs_reg_16_21_inst : DFF_X1 port map( D => N524, CK => clk, Q => n1972, QN 
                           => n26835);
   regs_nxt_reg_16_20_inst : DLH_X1 port map( G => n27580, D => n27282, Q => 
                           regs_nxt_16_20_port);
   regs_reg_16_20_inst : DFF_X1 port map( D => N523, CK => clk, Q => n1968, QN 
                           => n26834);
   regs_nxt_reg_16_19_inst : DLH_X1 port map( G => n27580, D => n27288, Q => 
                           regs_nxt_16_19_port);
   regs_reg_16_19_inst : DFF_X1 port map( D => N522, CK => clk, Q => n1964, QN 
                           => n26833);
   regs_nxt_reg_16_18_inst : DLH_X1 port map( G => n27582, D => n27294, Q => 
                           regs_nxt_16_18_port);
   regs_reg_16_18_inst : DFF_X1 port map( D => N521, CK => clk, Q => n1960, QN 
                           => n26832);
   regs_nxt_reg_16_17_inst : DLH_X1 port map( G => n27580, D => n27300, Q => 
                           regs_nxt_16_17_port);
   regs_reg_16_17_inst : DFF_X1 port map( D => N520, CK => clk, Q => n1956, QN 
                           => n26831);
   regs_nxt_reg_16_16_inst : DLH_X1 port map( G => n27582, D => n27306, Q => 
                           regs_nxt_16_16_port);
   regs_reg_16_16_inst : DFF_X1 port map( D => N519, CK => clk, Q => n1952, QN 
                           => n26830);
   regs_nxt_reg_16_15_inst : DLH_X1 port map( G => n27580, D => n27312, Q => 
                           regs_nxt_16_15_port);
   regs_reg_16_15_inst : DFF_X1 port map( D => N518, CK => clk, Q => n1948, QN 
                           => n26829);
   regs_nxt_reg_16_14_inst : DLH_X1 port map( G => n27582, D => n27318, Q => 
                           regs_nxt_16_14_port);
   regs_reg_16_14_inst : DFF_X1 port map( D => N517, CK => clk, Q => n1944, QN 
                           => n26828);
   regs_nxt_reg_16_13_inst : DLH_X1 port map( G => n27582, D => n27324, Q => 
                           regs_nxt_16_13_port);
   regs_reg_16_13_inst : DFF_X1 port map( D => N516, CK => clk, Q => n1940, QN 
                           => n26827);
   regs_nxt_reg_16_12_inst : DLH_X1 port map( G => n27582, D => n27330, Q => 
                           regs_nxt_16_12_port);
   regs_reg_16_12_inst : DFF_X1 port map( D => N515, CK => clk, Q => n1936, QN 
                           => n26826);
   regs_nxt_reg_16_11_inst : DLH_X1 port map( G => n27580, D => n27336, Q => 
                           regs_nxt_16_11_port);
   regs_reg_16_11_inst : DFF_X1 port map( D => N514, CK => clk, Q => n1932, QN 
                           => n26825);
   regs_nxt_reg_16_10_inst : DLH_X1 port map( G => n27580, D => n27342, Q => 
                           regs_nxt_16_10_port);
   regs_reg_16_10_inst : DFF_X1 port map( D => N513, CK => clk, Q => n1928, QN 
                           => n26824);
   regs_nxt_reg_16_9_inst : DLH_X1 port map( G => n27581, D => n27348, Q => 
                           regs_nxt_16_9_port);
   regs_reg_16_9_inst : DFF_X1 port map( D => N512, CK => clk, Q => n1924, QN 
                           => n26823);
   regs_nxt_reg_16_8_inst : DLH_X1 port map( G => n27581, D => n27354, Q => 
                           regs_nxt_16_8_port);
   regs_reg_16_8_inst : DFF_X1 port map( D => N511, CK => clk, Q => n1920, QN 
                           => n26822);
   regs_nxt_reg_16_7_inst : DLH_X1 port map( G => n27581, D => n27360, Q => 
                           regs_nxt_16_7_port);
   regs_reg_16_7_inst : DFF_X1 port map( D => N510, CK => clk, Q => n1916, QN 
                           => n26821);
   regs_nxt_reg_16_6_inst : DLH_X1 port map( G => n27581, D => n27366, Q => 
                           regs_nxt_16_6_port);
   regs_reg_16_6_inst : DFF_X1 port map( D => N509, CK => clk, Q => n1912, QN 
                           => n26820);
   regs_nxt_reg_16_5_inst : DLH_X1 port map( G => n27581, D => n27276, Q => 
                           regs_nxt_16_5_port);
   regs_reg_16_5_inst : DFF_X1 port map( D => N508, CK => clk, Q => n1908, QN 
                           => n26819);
   regs_nxt_reg_16_4_inst : DLH_X1 port map( G => n27581, D => n27438, Q => 
                           regs_nxt_16_4_port);
   regs_reg_16_4_inst : DFF_X1 port map( D => N507, CK => clk, Q => n1904, QN 
                           => n26818);
   regs_nxt_reg_16_3_inst : DLH_X1 port map( G => n27582, D => n27444, Q => 
                           regs_nxt_16_3_port);
   regs_reg_16_3_inst : DFF_X1 port map( D => N506, CK => clk, Q => n1900, QN 
                           => n26817);
   regs_nxt_reg_16_2_inst : DLH_X1 port map( G => n27581, D => n27450, Q => 
                           regs_nxt_16_2_port);
   regs_reg_16_2_inst : DFF_X1 port map( D => N505, CK => clk, Q => n1896, QN 
                           => n26816);
   regs_nxt_reg_16_1_inst : DLH_X1 port map( G => n27580, D => n27456, Q => 
                           regs_nxt_16_1_port);
   regs_reg_16_1_inst : DFF_X1 port map( D => N504, CK => clk, Q => n1892, QN 
                           => n26815);
   regs_nxt_reg_16_0_inst : DLH_X1 port map( G => n27581, D => n27464, Q => 
                           regs_nxt_16_0_port);
   regs_reg_16_0_inst : DFF_X1 port map( D => N503, CK => clk, Q => n1888, QN 
                           => n26814);
   regs_nxt_reg_17_31_inst : DLH_X1 port map( G => n27588, D => n27372, Q => 
                           regs_nxt_17_31_port);
   regs_reg_17_31_inst : DFF_X1 port map( D => N502, CK => clk, Q => n2610, QN 
                           => n26906);
   regs_nxt_reg_17_30_inst : DLH_X1 port map( G => n27588, D => n27378, Q => 
                           regs_nxt_17_30_port);
   regs_reg_17_30_inst : DFF_X1 port map( D => N501, CK => clk, Q => n2606, QN 
                           => n26905);
   regs_nxt_reg_17_29_inst : DLH_X1 port map( G => n27587, D => n27384, Q => 
                           regs_nxt_17_29_port);
   regs_reg_17_29_inst : DFF_X1 port map( D => N500, CK => clk, Q => n2602, QN 
                           => n26904);
   regs_nxt_reg_17_28_inst : DLH_X1 port map( G => n27587, D => n27390, Q => 
                           regs_nxt_17_28_port);
   regs_reg_17_28_inst : DFF_X1 port map( D => N499, CK => clk, Q => n2598, QN 
                           => n26903);
   regs_nxt_reg_17_27_inst : DLH_X1 port map( G => n27590, D => n27396, Q => 
                           regs_nxt_17_27_port);
   regs_reg_17_27_inst : DFF_X1 port map( D => N498, CK => clk, Q => n2594, QN 
                           => n26902);
   regs_nxt_reg_17_26_inst : DLH_X1 port map( G => n27589, D => n27402, Q => 
                           regs_nxt_17_26_port);
   regs_reg_17_26_inst : DFF_X1 port map( D => N497, CK => clk, Q => n2590, QN 
                           => n26901);
   regs_nxt_reg_17_25_inst : DLH_X1 port map( G => n27590, D => n27408, Q => 
                           regs_nxt_17_25_port);
   regs_reg_17_25_inst : DFF_X1 port map( D => N496, CK => clk, Q => n2586, QN 
                           => n26900);
   regs_nxt_reg_17_24_inst : DLH_X1 port map( G => n27589, D => n27414, Q => 
                           regs_nxt_17_24_port);
   regs_reg_17_24_inst : DFF_X1 port map( D => N495, CK => clk, Q => n2582, QN 
                           => n26899);
   regs_nxt_reg_17_23_inst : DLH_X1 port map( G => n27589, D => n27420, Q => 
                           regs_nxt_17_23_port);
   regs_reg_17_23_inst : DFF_X1 port map( D => N494, CK => clk, Q => n2578, QN 
                           => n26898);
   regs_nxt_reg_17_22_inst : DLH_X1 port map( G => n27589, D => n27426, Q => 
                           regs_nxt_17_22_port);
   regs_reg_17_22_inst : DFF_X1 port map( D => N493, CK => clk, Q => n2574, QN 
                           => n26897);
   regs_nxt_reg_17_21_inst : DLH_X1 port map( G => n27587, D => n27432, Q => 
                           regs_nxt_17_21_port);
   regs_reg_17_21_inst : DFF_X1 port map( D => N492, CK => clk, Q => n2570, QN 
                           => n26896);
   regs_nxt_reg_17_20_inst : DLH_X1 port map( G => n27587, D => n27282, Q => 
                           regs_nxt_17_20_port);
   regs_reg_17_20_inst : DFF_X1 port map( D => N491, CK => clk, Q => n2566, QN 
                           => n26895);
   regs_nxt_reg_17_19_inst : DLH_X1 port map( G => n27587, D => n27288, Q => 
                           regs_nxt_17_19_port);
   regs_reg_17_19_inst : DFF_X1 port map( D => N490, CK => clk, Q => n2562, QN 
                           => n26894);
   regs_nxt_reg_17_18_inst : DLH_X1 port map( G => n27589, D => n27294, Q => 
                           regs_nxt_17_18_port);
   regs_reg_17_18_inst : DFF_X1 port map( D => N489, CK => clk, Q => n2558, QN 
                           => n26893);
   regs_nxt_reg_17_17_inst : DLH_X1 port map( G => n27587, D => n27300, Q => 
                           regs_nxt_17_17_port);
   regs_reg_17_17_inst : DFF_X1 port map( D => N488, CK => clk, Q => n2554, QN 
                           => n26892);
   regs_nxt_reg_17_16_inst : DLH_X1 port map( G => n27589, D => n27306, Q => 
                           regs_nxt_17_16_port);
   regs_reg_17_16_inst : DFF_X1 port map( D => N487, CK => clk, Q => n2550, QN 
                           => n26891);
   regs_nxt_reg_17_15_inst : DLH_X1 port map( G => n27587, D => n27312, Q => 
                           regs_nxt_17_15_port);
   regs_reg_17_15_inst : DFF_X1 port map( D => N486, CK => clk, Q => n2546, QN 
                           => n26890);
   regs_nxt_reg_17_14_inst : DLH_X1 port map( G => n27589, D => n27318, Q => 
                           regs_nxt_17_14_port);
   regs_reg_17_14_inst : DFF_X1 port map( D => N485, CK => clk, Q => n_1439, QN
                           => n26599);
   regs_nxt_reg_17_13_inst : DLH_X1 port map( G => n27589, D => n27324, Q => 
                           regs_nxt_17_13_port);
   regs_reg_17_13_inst : DFF_X1 port map( D => N484, CK => clk, Q => n_1440, QN
                           => n26598);
   regs_nxt_reg_17_12_inst : DLH_X1 port map( G => n27589, D => n27330, Q => 
                           regs_nxt_17_12_port);
   regs_reg_17_12_inst : DFF_X1 port map( D => N483, CK => clk, Q => n_1441, QN
                           => n26597);
   regs_nxt_reg_17_11_inst : DLH_X1 port map( G => n27587, D => n27336, Q => 
                           regs_nxt_17_11_port);
   regs_reg_17_11_inst : DFF_X1 port map( D => N482, CK => clk, Q => n_1442, QN
                           => n26596);
   regs_nxt_reg_17_10_inst : DLH_X1 port map( G => n27587, D => n27342, Q => 
                           regs_nxt_17_10_port);
   regs_reg_17_10_inst : DFF_X1 port map( D => N481, CK => clk, Q => n_1443, QN
                           => n25269);
   regs_nxt_reg_17_9_inst : DLH_X1 port map( G => n27588, D => n27348, Q => 
                           regs_nxt_17_9_port);
   regs_reg_17_9_inst : DFF_X1 port map( D => N480, CK => clk, Q => n_1444, QN 
                           => n25268);
   regs_nxt_reg_17_8_inst : DLH_X1 port map( G => n27588, D => n27354, Q => 
                           regs_nxt_17_8_port);
   regs_reg_17_8_inst : DFF_X1 port map( D => N479, CK => clk, Q => n_1445, QN 
                           => n25267);
   regs_nxt_reg_17_7_inst : DLH_X1 port map( G => n27588, D => n27360, Q => 
                           regs_nxt_17_7_port);
   regs_reg_17_7_inst : DFF_X1 port map( D => N478, CK => clk, Q => n_1446, QN 
                           => n25266);
   regs_nxt_reg_17_6_inst : DLH_X1 port map( G => n27588, D => n27366, Q => 
                           regs_nxt_17_6_port);
   regs_reg_17_6_inst : DFF_X1 port map( D => N477, CK => clk, Q => n_1447, QN 
                           => n25265);
   regs_nxt_reg_17_5_inst : DLH_X1 port map( G => n27588, D => n27276, Q => 
                           regs_nxt_17_5_port);
   regs_reg_17_5_inst : DFF_X1 port map( D => N476, CK => clk, Q => n_1448, QN 
                           => n25264);
   regs_nxt_reg_17_4_inst : DLH_X1 port map( G => n27588, D => n27438, Q => 
                           regs_nxt_17_4_port);
   regs_reg_17_4_inst : DFF_X1 port map( D => N475, CK => clk, Q => n_1449, QN 
                           => n25263);
   regs_nxt_reg_17_3_inst : DLH_X1 port map( G => n27589, D => n27446, Q => 
                           regs_nxt_17_3_port);
   regs_reg_17_3_inst : DFF_X1 port map( D => N474, CK => clk, Q => n_1450, QN 
                           => n25262);
   regs_nxt_reg_17_2_inst : DLH_X1 port map( G => n27588, D => n27452, Q => 
                           regs_nxt_17_2_port);
   regs_reg_17_2_inst : DFF_X1 port map( D => N473, CK => clk, Q => n_1451, QN 
                           => n25261);
   regs_nxt_reg_17_1_inst : DLH_X1 port map( G => n27587, D => n27456, Q => 
                           regs_nxt_17_1_port);
   regs_reg_17_1_inst : DFF_X1 port map( D => N472, CK => clk, Q => n_1452, QN 
                           => n25260);
   regs_nxt_reg_17_0_inst : DLH_X1 port map( G => n27588, D => n27462, Q => 
                           regs_nxt_17_0_port);
   regs_reg_17_0_inst : DFF_X1 port map( D => N471, CK => clk, Q => n_1453, QN 
                           => n25259);
   regs_nxt_reg_18_31_inst : DLH_X1 port map( G => n27595, D => n27374, Q => 
                           regs_nxt_18_31_port);
   regs_reg_18_31_inst : DFF_X1 port map( D => N470, CK => clk, Q => 
                           regs_18_31_port, QN => n26961);
   regs_nxt_reg_18_30_inst : DLH_X1 port map( G => n27595, D => n27380, Q => 
                           regs_nxt_18_30_port);
   regs_reg_18_30_inst : DFF_X1 port map( D => N469, CK => clk, Q => 
                           regs_18_30_port, QN => n26960);
   regs_nxt_reg_18_29_inst : DLH_X1 port map( G => n27594, D => n27386, Q => 
                           regs_nxt_18_29_port);
   regs_reg_18_29_inst : DFF_X1 port map( D => N468, CK => clk, Q => 
                           regs_18_29_port, QN => n26959);
   regs_nxt_reg_18_28_inst : DLH_X1 port map( G => n27594, D => n27392, Q => 
                           regs_nxt_18_28_port);
   regs_reg_18_28_inst : DFF_X1 port map( D => N467, CK => clk, Q => 
                           regs_18_28_port, QN => n26958);
   regs_nxt_reg_18_27_inst : DLH_X1 port map( G => n27597, D => n27398, Q => 
                           regs_nxt_18_27_port);
   regs_reg_18_27_inst : DFF_X1 port map( D => N466, CK => clk, Q => 
                           regs_18_27_port, QN => n26957);
   regs_nxt_reg_18_26_inst : DLH_X1 port map( G => n27596, D => n27404, Q => 
                           regs_nxt_18_26_port);
   regs_reg_18_26_inst : DFF_X1 port map( D => N465, CK => clk, Q => 
                           regs_18_26_port, QN => n26956);
   regs_nxt_reg_18_25_inst : DLH_X1 port map( G => n27597, D => n27410, Q => 
                           regs_nxt_18_25_port);
   regs_reg_18_25_inst : DFF_X1 port map( D => N464, CK => clk, Q => 
                           regs_18_25_port, QN => n26955);
   regs_nxt_reg_18_24_inst : DLH_X1 port map( G => n27596, D => n27416, Q => 
                           regs_nxt_18_24_port);
   regs_reg_18_24_inst : DFF_X1 port map( D => N463, CK => clk, Q => 
                           regs_18_24_port, QN => n26954);
   regs_nxt_reg_18_23_inst : DLH_X1 port map( G => n27596, D => n27422, Q => 
                           regs_nxt_18_23_port);
   regs_reg_18_23_inst : DFF_X1 port map( D => N462, CK => clk, Q => 
                           regs_18_23_port, QN => n26953);
   regs_nxt_reg_18_22_inst : DLH_X1 port map( G => n27596, D => n27428, Q => 
                           regs_nxt_18_22_port);
   regs_reg_18_22_inst : DFF_X1 port map( D => N461, CK => clk, Q => 
                           regs_18_22_port, QN => n26952);
   regs_nxt_reg_18_21_inst : DLH_X1 port map( G => n27594, D => n27434, Q => 
                           regs_nxt_18_21_port);
   regs_reg_18_21_inst : DFF_X1 port map( D => N460, CK => clk, Q => 
                           regs_18_21_port, QN => n26951);
   regs_nxt_reg_18_20_inst : DLH_X1 port map( G => n27594, D => n27284, Q => 
                           regs_nxt_18_20_port);
   regs_reg_18_20_inst : DFF_X1 port map( D => N459, CK => clk, Q => 
                           regs_18_20_port, QN => n26950);
   regs_nxt_reg_18_19_inst : DLH_X1 port map( G => n27594, D => n27290, Q => 
                           regs_nxt_18_19_port);
   regs_reg_18_19_inst : DFF_X1 port map( D => N458, CK => clk, Q => 
                           regs_18_19_port, QN => n26949);
   regs_nxt_reg_18_18_inst : DLH_X1 port map( G => n27596, D => n27296, Q => 
                           regs_nxt_18_18_port);
   regs_reg_18_18_inst : DFF_X1 port map( D => N457, CK => clk, Q => 
                           regs_18_18_port, QN => n26948);
   regs_nxt_reg_18_17_inst : DLH_X1 port map( G => n27594, D => n27302, Q => 
                           regs_nxt_18_17_port);
   regs_reg_18_17_inst : DFF_X1 port map( D => N456, CK => clk, Q => 
                           regs_18_17_port, QN => n26947);
   regs_nxt_reg_18_16_inst : DLH_X1 port map( G => n27596, D => n27308, Q => 
                           regs_nxt_18_16_port);
   regs_reg_18_16_inst : DFF_X1 port map( D => N455, CK => clk, Q => 
                           regs_18_16_port, QN => n26946);
   regs_nxt_reg_18_15_inst : DLH_X1 port map( G => n27594, D => n27314, Q => 
                           regs_nxt_18_15_port);
   regs_reg_18_15_inst : DFF_X1 port map( D => N454, CK => clk, Q => 
                           regs_18_15_port, QN => n26945);
   regs_nxt_reg_18_14_inst : DLH_X1 port map( G => n27596, D => n27320, Q => 
                           regs_nxt_18_14_port);
   regs_reg_18_14_inst : DFF_X1 port map( D => N453, CK => clk, Q => 
                           regs_18_14_port, QN => n26944);
   regs_nxt_reg_18_13_inst : DLH_X1 port map( G => n27596, D => n27326, Q => 
                           regs_nxt_18_13_port);
   regs_reg_18_13_inst : DFF_X1 port map( D => N452, CK => clk, Q => 
                           regs_18_13_port, QN => n26943);
   regs_nxt_reg_18_12_inst : DLH_X1 port map( G => n27596, D => n27332, Q => 
                           regs_nxt_18_12_port);
   regs_reg_18_12_inst : DFF_X1 port map( D => N451, CK => clk, Q => 
                           regs_18_12_port, QN => n26942);
   regs_nxt_reg_18_11_inst : DLH_X1 port map( G => n27594, D => n27338, Q => 
                           regs_nxt_18_11_port);
   regs_reg_18_11_inst : DFF_X1 port map( D => N450, CK => clk, Q => 
                           regs_18_11_port, QN => n26941);
   regs_nxt_reg_18_10_inst : DLH_X1 port map( G => n27594, D => n27344, Q => 
                           regs_nxt_18_10_port);
   regs_reg_18_10_inst : DFF_X1 port map( D => N449, CK => clk, Q => 
                           regs_18_10_port, QN => n26940);
   regs_nxt_reg_18_9_inst : DLH_X1 port map( G => n27595, D => n27350, Q => 
                           regs_nxt_18_9_port);
   regs_reg_18_9_inst : DFF_X1 port map( D => N448, CK => clk, Q => 
                           regs_18_9_port, QN => n26939);
   regs_nxt_reg_18_8_inst : DLH_X1 port map( G => n27595, D => n27354, Q => 
                           regs_nxt_18_8_port);
   regs_reg_18_8_inst : DFF_X1 port map( D => N447, CK => clk, Q => 
                           regs_18_8_port, QN => n26938);
   regs_nxt_reg_18_7_inst : DLH_X1 port map( G => n27595, D => n27362, Q => 
                           regs_nxt_18_7_port);
   regs_reg_18_7_inst : DFF_X1 port map( D => N446, CK => clk, Q => 
                           regs_18_7_port, QN => n26937);
   regs_nxt_reg_18_6_inst : DLH_X1 port map( G => n27595, D => n27368, Q => 
                           regs_nxt_18_6_port);
   regs_reg_18_6_inst : DFF_X1 port map( D => N445, CK => clk, Q => 
                           regs_18_6_port, QN => n26936);
   regs_nxt_reg_18_5_inst : DLH_X1 port map( G => n27595, D => n27278, Q => 
                           regs_nxt_18_5_port);
   regs_reg_18_5_inst : DFF_X1 port map( D => N444, CK => clk, Q => 
                           regs_18_5_port, QN => n26935);
   regs_nxt_reg_18_4_inst : DLH_X1 port map( G => n27595, D => n27440, Q => 
                           regs_nxt_18_4_port);
   regs_reg_18_4_inst : DFF_X1 port map( D => N443, CK => clk, Q => 
                           regs_18_4_port, QN => n26934);
   regs_nxt_reg_18_3_inst : DLH_X1 port map( G => n27596, D => n27446, Q => 
                           regs_nxt_18_3_port);
   regs_reg_18_3_inst : DFF_X1 port map( D => N442, CK => clk, Q => 
                           regs_18_3_port, QN => n26933);
   regs_nxt_reg_18_2_inst : DLH_X1 port map( G => n27595, D => n27452, Q => 
                           regs_nxt_18_2_port);
   regs_reg_18_2_inst : DFF_X1 port map( D => N441, CK => clk, Q => 
                           regs_18_2_port, QN => n26932);
   regs_nxt_reg_18_1_inst : DLH_X1 port map( G => n27594, D => n27458, Q => 
                           regs_nxt_18_1_port);
   regs_reg_18_1_inst : DFF_X1 port map( D => N440, CK => clk, Q => 
                           regs_18_1_port, QN => n26931);
   regs_nxt_reg_18_0_inst : DLH_X1 port map( G => n27595, D => n27462, Q => 
                           regs_nxt_18_0_port);
   regs_reg_18_0_inst : DFF_X1 port map( D => N439, CK => clk, Q => 
                           regs_18_0_port, QN => n26930);
   regs_nxt_reg_19_31_inst : DLH_X1 port map( G => n27602, D => n27372, Q => 
                           regs_nxt_19_31_port);
   regs_reg_19_31_inst : DFF_X1 port map( D => N438, CK => clk, Q => n26442, QN
                           => n2611);
   regs_nxt_reg_19_30_inst : DLH_X1 port map( G => n27602, D => n27378, Q => 
                           regs_nxt_19_30_port);
   regs_reg_19_30_inst : DFF_X1 port map( D => N437, CK => clk, Q => n26441, QN
                           => n2607);
   regs_nxt_reg_19_29_inst : DLH_X1 port map( G => n27601, D => n27384, Q => 
                           regs_nxt_19_29_port);
   regs_reg_19_29_inst : DFF_X1 port map( D => N436, CK => clk, Q => n26440, QN
                           => n2603);
   regs_nxt_reg_19_28_inst : DLH_X1 port map( G => n27601, D => n27390, Q => 
                           regs_nxt_19_28_port);
   regs_reg_19_28_inst : DFF_X1 port map( D => N435, CK => clk, Q => n26439, QN
                           => n2599);
   regs_nxt_reg_19_27_inst : DLH_X1 port map( G => n27604, D => n27396, Q => 
                           regs_nxt_19_27_port);
   regs_reg_19_27_inst : DFF_X1 port map( D => N434, CK => clk, Q => n26438, QN
                           => n2595);
   regs_nxt_reg_19_26_inst : DLH_X1 port map( G => n27603, D => n27402, Q => 
                           regs_nxt_19_26_port);
   regs_reg_19_26_inst : DFF_X1 port map( D => N433, CK => clk, Q => n26437, QN
                           => n2591);
   regs_nxt_reg_19_25_inst : DLH_X1 port map( G => n27604, D => n27408, Q => 
                           regs_nxt_19_25_port);
   regs_reg_19_25_inst : DFF_X1 port map( D => N432, CK => clk, Q => n26436, QN
                           => n2587);
   regs_nxt_reg_19_24_inst : DLH_X1 port map( G => n27603, D => n27414, Q => 
                           regs_nxt_19_24_port);
   regs_reg_19_24_inst : DFF_X1 port map( D => N431, CK => clk, Q => n26435, QN
                           => n2583_port);
   regs_nxt_reg_19_23_inst : DLH_X1 port map( G => n27603, D => n27420, Q => 
                           regs_nxt_19_23_port);
   regs_reg_19_23_inst : DFF_X1 port map( D => N430, CK => clk, Q => n26434, QN
                           => n2579);
   regs_nxt_reg_19_22_inst : DLH_X1 port map( G => n27603, D => n27426, Q => 
                           regs_nxt_19_22_port);
   regs_reg_19_22_inst : DFF_X1 port map( D => N429, CK => clk, Q => n26433, QN
                           => n2575);
   regs_nxt_reg_19_21_inst : DLH_X1 port map( G => n27601, D => n27432, Q => 
                           regs_nxt_19_21_port);
   regs_reg_19_21_inst : DFF_X1 port map( D => N428, CK => clk, Q => n26432, QN
                           => n2571);
   regs_nxt_reg_19_20_inst : DLH_X1 port map( G => n27601, D => n27282, Q => 
                           regs_nxt_19_20_port);
   regs_reg_19_20_inst : DFF_X1 port map( D => N427, CK => clk, Q => n26431, QN
                           => n2567);
   regs_nxt_reg_19_19_inst : DLH_X1 port map( G => n27601, D => n27288, Q => 
                           regs_nxt_19_19_port);
   regs_reg_19_19_inst : DFF_X1 port map( D => N426, CK => clk, Q => n26430, QN
                           => n2563);
   regs_nxt_reg_19_18_inst : DLH_X1 port map( G => n27603, D => n27294, Q => 
                           regs_nxt_19_18_port);
   regs_reg_19_18_inst : DFF_X1 port map( D => N425, CK => clk, Q => n26429, QN
                           => n2559);
   regs_nxt_reg_19_17_inst : DLH_X1 port map( G => n27601, D => n27300, Q => 
                           regs_nxt_19_17_port);
   regs_reg_19_17_inst : DFF_X1 port map( D => N424, CK => clk, Q => n26428, QN
                           => n2555);
   regs_nxt_reg_19_16_inst : DLH_X1 port map( G => n27603, D => n27306, Q => 
                           regs_nxt_19_16_port);
   regs_reg_19_16_inst : DFF_X1 port map( D => N423, CK => clk, Q => n26427, QN
                           => n2551_port);
   regs_nxt_reg_19_15_inst : DLH_X1 port map( G => n27601, D => n27312, Q => 
                           regs_nxt_19_15_port);
   regs_reg_19_15_inst : DFF_X1 port map( D => N422, CK => clk, Q => n26426, QN
                           => n2547);
   regs_nxt_reg_19_14_inst : DLH_X1 port map( G => n27603, D => n27318, Q => 
                           regs_nxt_19_14_port);
   regs_reg_19_14_inst : DFF_X1 port map( D => N421, CK => clk, Q => n25448, QN
                           => n_1454);
   regs_nxt_reg_19_13_inst : DLH_X1 port map( G => n27603, D => n27324, Q => 
                           regs_nxt_19_13_port);
   regs_reg_19_13_inst : DFF_X1 port map( D => N420, CK => clk, Q => n25447, QN
                           => n_1455);
   regs_nxt_reg_19_12_inst : DLH_X1 port map( G => n27603, D => n27330, Q => 
                           regs_nxt_19_12_port);
   regs_reg_19_12_inst : DFF_X1 port map( D => N419, CK => clk, Q => n25446, QN
                           => n_1456);
   regs_nxt_reg_19_11_inst : DLH_X1 port map( G => n27601, D => n27336, Q => 
                           regs_nxt_19_11_port);
   regs_reg_19_11_inst : DFF_X1 port map( D => N418, CK => clk, Q => n25445, QN
                           => n_1457);
   regs_nxt_reg_19_10_inst : DLH_X1 port map( G => n27601, D => n27342, Q => 
                           regs_nxt_19_10_port);
   regs_reg_19_10_inst : DFF_X1 port map( D => N417, CK => clk, Q => n25444, QN
                           => n_1458);
   regs_nxt_reg_19_9_inst : DLH_X1 port map( G => n27602, D => n27348, Q => 
                           regs_nxt_19_9_port);
   regs_reg_19_9_inst : DFF_X1 port map( D => N416, CK => clk, Q => n25443, QN 
                           => n_1459);
   regs_nxt_reg_19_8_inst : DLH_X1 port map( G => n27602, D => n27354, Q => 
                           regs_nxt_19_8_port);
   regs_reg_19_8_inst : DFF_X1 port map( D => N415, CK => clk, Q => n25442, QN 
                           => n_1460);
   regs_nxt_reg_19_7_inst : DLH_X1 port map( G => n27602, D => n27360, Q => 
                           regs_nxt_19_7_port);
   regs_reg_19_7_inst : DFF_X1 port map( D => N414, CK => clk, Q => n25441, QN 
                           => n_1461);
   regs_nxt_reg_19_6_inst : DLH_X1 port map( G => n27602, D => n27366, Q => 
                           regs_nxt_19_6_port);
   regs_reg_19_6_inst : DFF_X1 port map( D => N413, CK => clk, Q => n25440, QN 
                           => n_1462);
   regs_nxt_reg_19_5_inst : DLH_X1 port map( G => n27602, D => n27276, Q => 
                           regs_nxt_19_5_port);
   regs_reg_19_5_inst : DFF_X1 port map( D => N412, CK => clk, Q => n25439, QN 
                           => n_1463);
   regs_nxt_reg_19_4_inst : DLH_X1 port map( G => n27602, D => n27438, Q => 
                           regs_nxt_19_4_port);
   regs_reg_19_4_inst : DFF_X1 port map( D => N411, CK => clk, Q => n25438, QN 
                           => n_1464);
   regs_nxt_reg_19_3_inst : DLH_X1 port map( G => n27603, D => n27446, Q => 
                           regs_nxt_19_3_port);
   regs_reg_19_3_inst : DFF_X1 port map( D => N410, CK => clk, Q => n25437, QN 
                           => n_1465);
   regs_nxt_reg_19_2_inst : DLH_X1 port map( G => n27602, D => n27452, Q => 
                           regs_nxt_19_2_port);
   regs_reg_19_2_inst : DFF_X1 port map( D => N409, CK => clk, Q => n25436, QN 
                           => n_1466);
   regs_nxt_reg_19_1_inst : DLH_X1 port map( G => n27601, D => n27456, Q => 
                           regs_nxt_19_1_port);
   regs_reg_19_1_inst : DFF_X1 port map( D => N408, CK => clk, Q => n25435, QN 
                           => n_1467);
   regs_nxt_reg_19_0_inst : DLH_X1 port map( G => n27602, D => n27462, Q => 
                           regs_nxt_19_0_port);
   regs_reg_19_0_inst : DFF_X1 port map( D => N407, CK => clk, Q => n25434, QN 
                           => n_1468);
   regs_nxt_reg_20_31_inst : DLH_X1 port map( G => n27609, D => n27374, Q => 
                           regs_nxt_20_31_port);
   regs_reg_20_31_inst : DFF_X1 port map( D => N406, CK => clk, Q => n2609, QN 
                           => n26588);
   regs_nxt_reg_20_30_inst : DLH_X1 port map( G => n27609, D => n27380, Q => 
                           regs_nxt_20_30_port);
   regs_reg_20_30_inst : DFF_X1 port map( D => N405, CK => clk, Q => n2605, QN 
                           => n26587);
   regs_nxt_reg_20_29_inst : DLH_X1 port map( G => n27608, D => n27386, Q => 
                           regs_nxt_20_29_port);
   regs_reg_20_29_inst : DFF_X1 port map( D => N404, CK => clk, Q => n2601, QN 
                           => n26586);
   regs_nxt_reg_20_28_inst : DLH_X1 port map( G => n27608, D => n27392, Q => 
                           regs_nxt_20_28_port);
   regs_reg_20_28_inst : DFF_X1 port map( D => N403, CK => clk, Q => n2597, QN 
                           => n26585);
   regs_nxt_reg_20_27_inst : DLH_X1 port map( G => n27611, D => n27398, Q => 
                           regs_nxt_20_27_port);
   regs_reg_20_27_inst : DFF_X1 port map( D => N402, CK => clk, Q => n2593, QN 
                           => n26584);
   regs_nxt_reg_20_26_inst : DLH_X1 port map( G => n27610, D => n27404, Q => 
                           regs_nxt_20_26_port);
   regs_reg_20_26_inst : DFF_X1 port map( D => N401, CK => clk, Q => n2589, QN 
                           => n26583);
   regs_nxt_reg_20_25_inst : DLH_X1 port map( G => n27611, D => n27410, Q => 
                           regs_nxt_20_25_port);
   regs_reg_20_25_inst : DFF_X1 port map( D => N400, CK => clk, Q => n2585, QN 
                           => n26582);
   regs_nxt_reg_20_24_inst : DLH_X1 port map( G => n27610, D => n27416, Q => 
                           regs_nxt_20_24_port);
   regs_reg_20_24_inst : DFF_X1 port map( D => N399, CK => clk, Q => n2581, QN 
                           => n26581);
   regs_nxt_reg_20_23_inst : DLH_X1 port map( G => n27610, D => n27422, Q => 
                           regs_nxt_20_23_port);
   regs_reg_20_23_inst : DFF_X1 port map( D => N398, CK => clk, Q => n2577, QN 
                           => n26580);
   regs_nxt_reg_20_22_inst : DLH_X1 port map( G => n27610, D => n27428, Q => 
                           regs_nxt_20_22_port);
   regs_reg_20_22_inst : DFF_X1 port map( D => N397, CK => clk, Q => n2573, QN 
                           => n26579);
   regs_nxt_reg_20_21_inst : DLH_X1 port map( G => n27608, D => n27434, Q => 
                           regs_nxt_20_21_port);
   regs_reg_20_21_inst : DFF_X1 port map( D => N396, CK => clk, Q => n2569, QN 
                           => n26578);
   regs_nxt_reg_20_20_inst : DLH_X1 port map( G => n27608, D => n27284, Q => 
                           regs_nxt_20_20_port);
   regs_reg_20_20_inst : DFF_X1 port map( D => N395, CK => clk, Q => n2565, QN 
                           => n26577);
   regs_nxt_reg_20_19_inst : DLH_X1 port map( G => n27608, D => n27290, Q => 
                           regs_nxt_20_19_port);
   regs_reg_20_19_inst : DFF_X1 port map( D => N394, CK => clk, Q => n2561, QN 
                           => n26576);
   regs_nxt_reg_20_18_inst : DLH_X1 port map( G => n27610, D => n27296, Q => 
                           regs_nxt_20_18_port);
   regs_reg_20_18_inst : DFF_X1 port map( D => N393, CK => clk, Q => n2557, QN 
                           => n26575);
   regs_nxt_reg_20_17_inst : DLH_X1 port map( G => n27608, D => n27302, Q => 
                           regs_nxt_20_17_port);
   regs_reg_20_17_inst : DFF_X1 port map( D => N392, CK => clk, Q => n2553, QN 
                           => n26574);
   regs_nxt_reg_20_16_inst : DLH_X1 port map( G => n27610, D => n27308, Q => 
                           regs_nxt_20_16_port);
   regs_reg_20_16_inst : DFF_X1 port map( D => N391, CK => clk, Q => n26697, QN
                           => n25516);
   regs_nxt_reg_20_15_inst : DLH_X1 port map( G => n27608, D => n27314, Q => 
                           regs_nxt_20_15_port);
   regs_reg_20_15_inst : DFF_X1 port map( D => N390, CK => clk, Q => n26696, QN
                           => n25515);
   regs_nxt_reg_20_14_inst : DLH_X1 port map( G => n27610, D => n27320, Q => 
                           regs_nxt_20_14_port);
   regs_reg_20_14_inst : DFF_X1 port map( D => N389, CK => clk, Q => n_1469, QN
                           => n25514);
   regs_nxt_reg_20_13_inst : DLH_X1 port map( G => n27610, D => n27326, Q => 
                           regs_nxt_20_13_port);
   regs_reg_20_13_inst : DFF_X1 port map( D => N388, CK => clk, Q => n_1470, QN
                           => n25513);
   regs_nxt_reg_20_12_inst : DLH_X1 port map( G => n27610, D => n27332, Q => 
                           regs_nxt_20_12_port);
   regs_reg_20_12_inst : DFF_X1 port map( D => N387, CK => clk, Q => n_1471, QN
                           => n25512);
   regs_nxt_reg_20_11_inst : DLH_X1 port map( G => n27608, D => n27338, Q => 
                           regs_nxt_20_11_port);
   regs_reg_20_11_inst : DFF_X1 port map( D => N386, CK => clk, Q => n_1472, QN
                           => n25511);
   regs_nxt_reg_20_10_inst : DLH_X1 port map( G => n27608, D => n27344, Q => 
                           regs_nxt_20_10_port);
   regs_reg_20_10_inst : DFF_X1 port map( D => N385, CK => clk, Q => n_1473, QN
                           => n25510);
   regs_nxt_reg_20_9_inst : DLH_X1 port map( G => n27609, D => n27350, Q => 
                           regs_nxt_20_9_port);
   regs_reg_20_9_inst : DFF_X1 port map( D => N384, CK => clk, Q => n_1474, QN 
                           => n25509);
   regs_nxt_reg_20_8_inst : DLH_X1 port map( G => n27609, D => n27356, Q => 
                           regs_nxt_20_8_port);
   regs_reg_20_8_inst : DFF_X1 port map( D => N383, CK => clk, Q => n_1475, QN 
                           => n25508);
   regs_nxt_reg_20_7_inst : DLH_X1 port map( G => n27609, D => n27362, Q => 
                           regs_nxt_20_7_port);
   regs_reg_20_7_inst : DFF_X1 port map( D => N382, CK => clk, Q => n_1476, QN 
                           => n25507);
   regs_nxt_reg_20_6_inst : DLH_X1 port map( G => n27609, D => n27368, Q => 
                           regs_nxt_20_6_port);
   regs_reg_20_6_inst : DFF_X1 port map( D => N381, CK => clk, Q => n_1477, QN 
                           => n25506);
   regs_nxt_reg_20_5_inst : DLH_X1 port map( G => n27609, D => n27278, Q => 
                           regs_nxt_20_5_port);
   regs_reg_20_5_inst : DFF_X1 port map( D => N380, CK => clk, Q => n_1478, QN 
                           => n25505);
   regs_nxt_reg_20_4_inst : DLH_X1 port map( G => n27609, D => n27440, Q => 
                           regs_nxt_20_4_port);
   regs_reg_20_4_inst : DFF_X1 port map( D => N379, CK => clk, Q => n_1479, QN 
                           => n25504);
   regs_nxt_reg_20_3_inst : DLH_X1 port map( G => n27610, D => n27446, Q => 
                           regs_nxt_20_3_port);
   regs_reg_20_3_inst : DFF_X1 port map( D => N378, CK => clk, Q => n_1480, QN 
                           => n25503);
   regs_nxt_reg_20_2_inst : DLH_X1 port map( G => n27609, D => n27452, Q => 
                           regs_nxt_20_2_port);
   regs_reg_20_2_inst : DFF_X1 port map( D => N377, CK => clk, Q => n_1481, QN 
                           => n25502);
   regs_nxt_reg_20_1_inst : DLH_X1 port map( G => n27608, D => n27458, Q => 
                           regs_nxt_20_1_port);
   regs_reg_20_1_inst : DFF_X1 port map( D => N376, CK => clk, Q => n_1482, QN 
                           => n25501);
   regs_nxt_reg_20_0_inst : DLH_X1 port map( G => n27609, D => n27464, Q => 
                           regs_nxt_20_0_port);
   regs_reg_20_0_inst : DFF_X1 port map( D => N375, CK => clk, Q => n_1483, QN 
                           => n25500);
   regs_nxt_reg_21_31_inst : DLH_X1 port map( G => n27616, D => n27374, Q => 
                           regs_nxt_21_31_port);
   regs_reg_21_31_inst : DFF_X1 port map( D => N374, CK => clk, Q => n26813, QN
                           => n2014);
   regs_nxt_reg_21_30_inst : DLH_X1 port map( G => n27616, D => n27380, Q => 
                           regs_nxt_21_30_port);
   regs_reg_21_30_inst : DFF_X1 port map( D => N373, CK => clk, Q => n26812, QN
                           => n2010);
   regs_nxt_reg_21_29_inst : DLH_X1 port map( G => n27615, D => n27386, Q => 
                           regs_nxt_21_29_port);
   regs_reg_21_29_inst : DFF_X1 port map( D => N372, CK => clk, Q => n26811, QN
                           => n2006);
   regs_nxt_reg_21_28_inst : DLH_X1 port map( G => n27615, D => n27392, Q => 
                           regs_nxt_21_28_port);
   regs_reg_21_28_inst : DFF_X1 port map( D => N371, CK => clk, Q => n26810, QN
                           => n2002);
   regs_nxt_reg_21_27_inst : DLH_X1 port map( G => n27618, D => n27398, Q => 
                           regs_nxt_21_27_port);
   regs_reg_21_27_inst : DFF_X1 port map( D => N370, CK => clk, Q => n26809, QN
                           => n1998);
   regs_nxt_reg_21_26_inst : DLH_X1 port map( G => n27617, D => n27404, Q => 
                           regs_nxt_21_26_port);
   regs_reg_21_26_inst : DFF_X1 port map( D => N369, CK => clk, Q => n26808, QN
                           => n1994);
   regs_nxt_reg_21_25_inst : DLH_X1 port map( G => n27618, D => n27410, Q => 
                           regs_nxt_21_25_port);
   regs_reg_21_25_inst : DFF_X1 port map( D => N368, CK => clk, Q => n26807, QN
                           => n1990);
   regs_nxt_reg_21_24_inst : DLH_X1 port map( G => n27617, D => n27416, Q => 
                           regs_nxt_21_24_port);
   regs_reg_21_24_inst : DFF_X1 port map( D => N367, CK => clk, Q => n26806, QN
                           => n1986);
   regs_nxt_reg_21_23_inst : DLH_X1 port map( G => n27617, D => n27422, Q => 
                           regs_nxt_21_23_port);
   regs_reg_21_23_inst : DFF_X1 port map( D => N366, CK => clk, Q => n26805, QN
                           => n1982);
   regs_nxt_reg_21_22_inst : DLH_X1 port map( G => n27617, D => n27428, Q => 
                           regs_nxt_21_22_port);
   regs_reg_21_22_inst : DFF_X1 port map( D => N365, CK => clk, Q => n26804, QN
                           => n1978);
   regs_nxt_reg_21_21_inst : DLH_X1 port map( G => n27615, D => n27434, Q => 
                           regs_nxt_21_21_port);
   regs_reg_21_21_inst : DFF_X1 port map( D => N364, CK => clk, Q => n26803, QN
                           => n1974);
   regs_nxt_reg_21_20_inst : DLH_X1 port map( G => n27615, D => n27284, Q => 
                           regs_nxt_21_20_port);
   regs_reg_21_20_inst : DFF_X1 port map( D => N363, CK => clk, Q => n26802, QN
                           => n1970);
   regs_nxt_reg_21_19_inst : DLH_X1 port map( G => n27615, D => n27290, Q => 
                           regs_nxt_21_19_port);
   regs_reg_21_19_inst : DFF_X1 port map( D => N362, CK => clk, Q => n26801, QN
                           => n1966);
   regs_nxt_reg_21_18_inst : DLH_X1 port map( G => n27617, D => n27296, Q => 
                           regs_nxt_21_18_port);
   regs_reg_21_18_inst : DFF_X1 port map( D => N361, CK => clk, Q => n26800, QN
                           => n1962);
   regs_nxt_reg_21_17_inst : DLH_X1 port map( G => n27615, D => n27302, Q => 
                           regs_nxt_21_17_port);
   regs_reg_21_17_inst : DFF_X1 port map( D => N360, CK => clk, Q => n26799, QN
                           => n1958);
   regs_nxt_reg_21_16_inst : DLH_X1 port map( G => n27617, D => n27308, Q => 
                           regs_nxt_21_16_port);
   regs_reg_21_16_inst : DFF_X1 port map( D => N359, CK => clk, Q => n26798, QN
                           => n1954);
   regs_nxt_reg_21_15_inst : DLH_X1 port map( G => n27615, D => n27314, Q => 
                           regs_nxt_21_15_port);
   regs_reg_21_15_inst : DFF_X1 port map( D => N358, CK => clk, Q => n26797, QN
                           => n1950);
   regs_nxt_reg_21_14_inst : DLH_X1 port map( G => n27617, D => n27320, Q => 
                           regs_nxt_21_14_port);
   regs_reg_21_14_inst : DFF_X1 port map( D => N357, CK => clk, Q => n26796, QN
                           => n1946);
   regs_nxt_reg_21_13_inst : DLH_X1 port map( G => n27617, D => n27326, Q => 
                           regs_nxt_21_13_port);
   regs_reg_21_13_inst : DFF_X1 port map( D => N356, CK => clk, Q => n26795, QN
                           => n1942);
   regs_nxt_reg_21_12_inst : DLH_X1 port map( G => n27617, D => n27332, Q => 
                           regs_nxt_21_12_port);
   regs_reg_21_12_inst : DFF_X1 port map( D => N355, CK => clk, Q => n26794, QN
                           => n1938);
   regs_nxt_reg_21_11_inst : DLH_X1 port map( G => n27615, D => n27338, Q => 
                           regs_nxt_21_11_port);
   regs_reg_21_11_inst : DFF_X1 port map( D => N354, CK => clk, Q => n26793, QN
                           => n1934);
   regs_nxt_reg_21_10_inst : DLH_X1 port map( G => n27615, D => n27344, Q => 
                           regs_nxt_21_10_port);
   regs_reg_21_10_inst : DFF_X1 port map( D => N353, CK => clk, Q => n26792, QN
                           => n1930);
   regs_nxt_reg_21_9_inst : DLH_X1 port map( G => n27616, D => n27350, Q => 
                           regs_nxt_21_9_port);
   regs_reg_21_9_inst : DFF_X1 port map( D => N352, CK => clk, Q => n26791, QN 
                           => n1926);
   regs_nxt_reg_21_8_inst : DLH_X1 port map( G => n27616, D => n27356, Q => 
                           regs_nxt_21_8_port);
   regs_reg_21_8_inst : DFF_X1 port map( D => N351, CK => clk, Q => n26790, QN 
                           => n1922);
   regs_nxt_reg_21_7_inst : DLH_X1 port map( G => n27616, D => n27362, Q => 
                           regs_nxt_21_7_port);
   regs_reg_21_7_inst : DFF_X1 port map( D => N350, CK => clk, Q => n26789, QN 
                           => n1918);
   regs_nxt_reg_21_6_inst : DLH_X1 port map( G => n27616, D => n27368, Q => 
                           regs_nxt_21_6_port);
   regs_reg_21_6_inst : DFF_X1 port map( D => N349, CK => clk, Q => n26788, QN 
                           => n1914);
   regs_nxt_reg_21_5_inst : DLH_X1 port map( G => n27616, D => n27278, Q => 
                           regs_nxt_21_5_port);
   regs_reg_21_5_inst : DFF_X1 port map( D => N348, CK => clk, Q => n26787, QN 
                           => n1910);
   regs_nxt_reg_21_4_inst : DLH_X1 port map( G => n27616, D => n27440, Q => 
                           regs_nxt_21_4_port);
   regs_reg_21_4_inst : DFF_X1 port map( D => N347, CK => clk, Q => n26786, QN 
                           => n1906);
   regs_nxt_reg_21_3_inst : DLH_X1 port map( G => n27617, D => n27446, Q => 
                           regs_nxt_21_3_port);
   regs_reg_21_3_inst : DFF_X1 port map( D => N346, CK => clk, Q => n26785, QN 
                           => n1902);
   regs_nxt_reg_21_2_inst : DLH_X1 port map( G => n27616, D => n27452, Q => 
                           regs_nxt_21_2_port);
   regs_reg_21_2_inst : DFF_X1 port map( D => N345, CK => clk, Q => n26784, QN 
                           => n1898);
   regs_nxt_reg_21_1_inst : DLH_X1 port map( G => n27615, D => n27458, Q => 
                           regs_nxt_21_1_port);
   regs_reg_21_1_inst : DFF_X1 port map( D => N344, CK => clk, Q => n26783, QN 
                           => n1894);
   regs_nxt_reg_21_0_inst : DLH_X1 port map( G => n27616, D => n27464, Q => 
                           regs_nxt_21_0_port);
   regs_reg_21_0_inst : DFF_X1 port map( D => N343, CK => clk, Q => n26782, QN 
                           => n1890);
   regs_nxt_reg_22_31_inst : DLH_X1 port map( G => n27623, D => n27373, Q => 
                           regs_nxt_22_31_port);
   regs_reg_22_31_inst : DFF_X1 port map( D => N342, CK => clk, Q => n2011, QN 
                           => n26529);
   regs_nxt_reg_22_30_inst : DLH_X1 port map( G => n27623, D => n27379, Q => 
                           regs_nxt_22_30_port);
   regs_reg_22_30_inst : DFF_X1 port map( D => N341, CK => clk, Q => n2007, QN 
                           => n26528);
   regs_nxt_reg_22_29_inst : DLH_X1 port map( G => n27622, D => n27385, Q => 
                           regs_nxt_22_29_port);
   regs_reg_22_29_inst : DFF_X1 port map( D => N340, CK => clk, Q => n2003, QN 
                           => n26527);
   regs_nxt_reg_22_28_inst : DLH_X1 port map( G => n27622, D => n27391, Q => 
                           regs_nxt_22_28_port);
   regs_reg_22_28_inst : DFF_X1 port map( D => N339, CK => clk, Q => n1999, QN 
                           => n26526);
   regs_nxt_reg_22_27_inst : DLH_X1 port map( G => n27625, D => n27397, Q => 
                           regs_nxt_22_27_port);
   regs_reg_22_27_inst : DFF_X1 port map( D => N338, CK => clk, Q => n1995, QN 
                           => n26525);
   regs_nxt_reg_22_26_inst : DLH_X1 port map( G => n27624, D => n27403, Q => 
                           regs_nxt_22_26_port);
   regs_reg_22_26_inst : DFF_X1 port map( D => N337, CK => clk, Q => n1991, QN 
                           => n26524);
   regs_nxt_reg_22_25_inst : DLH_X1 port map( G => n27625, D => n27409, Q => 
                           regs_nxt_22_25_port);
   regs_reg_22_25_inst : DFF_X1 port map( D => N336, CK => clk, Q => n1987, QN 
                           => n26523);
   regs_nxt_reg_22_24_inst : DLH_X1 port map( G => n27624, D => n27415, Q => 
                           regs_nxt_22_24_port);
   regs_reg_22_24_inst : DFF_X1 port map( D => N335, CK => clk, Q => n1983, QN 
                           => n26522);
   regs_nxt_reg_22_23_inst : DLH_X1 port map( G => n27624, D => n27421, Q => 
                           regs_nxt_22_23_port);
   regs_reg_22_23_inst : DFF_X1 port map( D => N334, CK => clk, Q => n1979, QN 
                           => n26521);
   regs_nxt_reg_22_22_inst : DLH_X1 port map( G => n27624, D => n27427, Q => 
                           regs_nxt_22_22_port);
   regs_reg_22_22_inst : DFF_X1 port map( D => N333, CK => clk, Q => n1975, QN 
                           => n26520);
   regs_nxt_reg_22_21_inst : DLH_X1 port map( G => n27622, D => n27433, Q => 
                           regs_nxt_22_21_port);
   regs_reg_22_21_inst : DFF_X1 port map( D => N332, CK => clk, Q => n1971, QN 
                           => n26519);
   regs_nxt_reg_22_20_inst : DLH_X1 port map( G => n27622, D => n27283, Q => 
                           regs_nxt_22_20_port);
   regs_reg_22_20_inst : DFF_X1 port map( D => N331, CK => clk, Q => n1967, QN 
                           => n26518);
   regs_nxt_reg_22_19_inst : DLH_X1 port map( G => n27622, D => n27289, Q => 
                           regs_nxt_22_19_port);
   regs_reg_22_19_inst : DFF_X1 port map( D => N330, CK => clk, Q => n1963, QN 
                           => n26517);
   regs_nxt_reg_22_18_inst : DLH_X1 port map( G => n27624, D => n27295, Q => 
                           regs_nxt_22_18_port);
   regs_reg_22_18_inst : DFF_X1 port map( D => N329, CK => clk, Q => n1959, QN 
                           => n26516);
   regs_nxt_reg_22_17_inst : DLH_X1 port map( G => n27622, D => n27301, Q => 
                           regs_nxt_22_17_port);
   regs_reg_22_17_inst : DFF_X1 port map( D => N328, CK => clk, Q => n1955, QN 
                           => n26515);
   regs_nxt_reg_22_16_inst : DLH_X1 port map( G => n27624, D => n27307, Q => 
                           regs_nxt_22_16_port);
   regs_reg_22_16_inst : DFF_X1 port map( D => N327, CK => clk, Q => n1951, QN 
                           => n26514);
   regs_nxt_reg_22_15_inst : DLH_X1 port map( G => n27622, D => n27313, Q => 
                           regs_nxt_22_15_port);
   regs_reg_22_15_inst : DFF_X1 port map( D => N326, CK => clk, Q => n1947, QN 
                           => n26513);
   regs_nxt_reg_22_14_inst : DLH_X1 port map( G => n27624, D => n27319, Q => 
                           regs_nxt_22_14_port);
   regs_reg_22_14_inst : DFF_X1 port map( D => N325, CK => clk, Q => n1943, QN 
                           => n26512);
   regs_nxt_reg_22_13_inst : DLH_X1 port map( G => n27624, D => n27325, Q => 
                           regs_nxt_22_13_port);
   regs_reg_22_13_inst : DFF_X1 port map( D => N324, CK => clk, Q => n1939, QN 
                           => n26511);
   regs_nxt_reg_22_12_inst : DLH_X1 port map( G => n27624, D => n27331, Q => 
                           regs_nxt_22_12_port);
   regs_reg_22_12_inst : DFF_X1 port map( D => N323, CK => clk, Q => n1935, QN 
                           => n26510);
   regs_nxt_reg_22_11_inst : DLH_X1 port map( G => n27622, D => n27337, Q => 
                           regs_nxt_22_11_port);
   regs_reg_22_11_inst : DFF_X1 port map( D => N322, CK => clk, Q => n1931, QN 
                           => n26509);
   regs_nxt_reg_22_10_inst : DLH_X1 port map( G => n27622, D => n27343, Q => 
                           regs_nxt_22_10_port);
   regs_reg_22_10_inst : DFF_X1 port map( D => N321, CK => clk, Q => n1927, QN 
                           => n26508);
   regs_nxt_reg_22_9_inst : DLH_X1 port map( G => n27623, D => n27349, Q => 
                           regs_nxt_22_9_port);
   regs_reg_22_9_inst : DFF_X1 port map( D => N320, CK => clk, Q => n1923, QN 
                           => n26507);
   regs_nxt_reg_22_8_inst : DLH_X1 port map( G => n27623, D => n27356, Q => 
                           regs_nxt_22_8_port);
   regs_reg_22_8_inst : DFF_X1 port map( D => N319, CK => clk, Q => n1919, QN 
                           => n26506);
   regs_nxt_reg_22_7_inst : DLH_X1 port map( G => n27623, D => n27361, Q => 
                           regs_nxt_22_7_port);
   regs_reg_22_7_inst : DFF_X1 port map( D => N318, CK => clk, Q => n1915, QN 
                           => n26505);
   regs_nxt_reg_22_6_inst : DLH_X1 port map( G => n27623, D => n27367, Q => 
                           regs_nxt_22_6_port);
   regs_reg_22_6_inst : DFF_X1 port map( D => N317, CK => clk, Q => n1911, QN 
                           => n26504);
   regs_nxt_reg_22_5_inst : DLH_X1 port map( G => n27623, D => n27277, Q => 
                           regs_nxt_22_5_port);
   regs_reg_22_5_inst : DFF_X1 port map( D => N316, CK => clk, Q => n1907, QN 
                           => n26503);
   regs_nxt_reg_22_4_inst : DLH_X1 port map( G => n27623, D => n27439, Q => 
                           regs_nxt_22_4_port);
   regs_reg_22_4_inst : DFF_X1 port map( D => N315, CK => clk, Q => n1903, QN 
                           => n26502);
   regs_nxt_reg_22_3_inst : DLH_X1 port map( G => n27624, D => n27445, Q => 
                           regs_nxt_22_3_port);
   regs_reg_22_3_inst : DFF_X1 port map( D => N314, CK => clk, Q => n1899, QN 
                           => n26501);
   regs_nxt_reg_22_2_inst : DLH_X1 port map( G => n27623, D => n27451, Q => 
                           regs_nxt_22_2_port);
   regs_reg_22_2_inst : DFF_X1 port map( D => N313, CK => clk, Q => n1895, QN 
                           => n26500);
   regs_nxt_reg_22_1_inst : DLH_X1 port map( G => n27622, D => n27457, Q => 
                           regs_nxt_22_1_port);
   regs_reg_22_1_inst : DFF_X1 port map( D => N312, CK => clk, Q => n1891, QN 
                           => n26499);
   regs_nxt_reg_22_0_inst : DLH_X1 port map( G => n27623, D => n27463, Q => 
                           regs_nxt_22_0_port);
   regs_reg_22_0_inst : DFF_X1 port map( D => N311, CK => clk, Q => n1887, QN 
                           => n26498);
   regs_nxt_reg_23_31_inst : DLH_X1 port map( G => n27630, D => n27373, Q => 
                           regs_nxt_23_31_port);
   regs_reg_23_31_inst : DFF_X1 port map( D => N310, CK => clk, Q => n26474, QN
                           => n2013);
   regs_nxt_reg_23_30_inst : DLH_X1 port map( G => n27630, D => n27379, Q => 
                           regs_nxt_23_30_port);
   regs_reg_23_30_inst : DFF_X1 port map( D => N309, CK => clk, Q => n26473, QN
                           => n2009);
   regs_nxt_reg_23_29_inst : DLH_X1 port map( G => n27629, D => n27385, Q => 
                           regs_nxt_23_29_port);
   regs_reg_23_29_inst : DFF_X1 port map( D => N308, CK => clk, Q => n26472, QN
                           => n2005);
   regs_nxt_reg_23_28_inst : DLH_X1 port map( G => n27629, D => n27391, Q => 
                           regs_nxt_23_28_port);
   regs_reg_23_28_inst : DFF_X1 port map( D => N307, CK => clk, Q => n26471, QN
                           => n2001);
   regs_nxt_reg_23_27_inst : DLH_X1 port map( G => n27632, D => n27397, Q => 
                           regs_nxt_23_27_port);
   regs_reg_23_27_inst : DFF_X1 port map( D => N306, CK => clk, Q => n26470, QN
                           => n1997);
   regs_nxt_reg_23_26_inst : DLH_X1 port map( G => n27631, D => n27403, Q => 
                           regs_nxt_23_26_port);
   regs_reg_23_26_inst : DFF_X1 port map( D => N305, CK => clk, Q => n26469, QN
                           => n1993);
   regs_nxt_reg_23_25_inst : DLH_X1 port map( G => n27632, D => n27409, Q => 
                           regs_nxt_23_25_port);
   regs_reg_23_25_inst : DFF_X1 port map( D => N304, CK => clk, Q => n26468, QN
                           => n1989);
   regs_nxt_reg_23_24_inst : DLH_X1 port map( G => n27631, D => n27415, Q => 
                           regs_nxt_23_24_port);
   regs_reg_23_24_inst : DFF_X1 port map( D => N303, CK => clk, Q => n26467, QN
                           => n1985);
   regs_nxt_reg_23_23_inst : DLH_X1 port map( G => n27631, D => n27421, Q => 
                           regs_nxt_23_23_port);
   regs_reg_23_23_inst : DFF_X1 port map( D => N302, CK => clk, Q => n26466, QN
                           => n1981);
   regs_nxt_reg_23_22_inst : DLH_X1 port map( G => n27631, D => n27427, Q => 
                           regs_nxt_23_22_port);
   regs_reg_23_22_inst : DFF_X1 port map( D => N301, CK => clk, Q => n26465, QN
                           => n1977);
   regs_nxt_reg_23_21_inst : DLH_X1 port map( G => n27629, D => n27433, Q => 
                           regs_nxt_23_21_port);
   regs_reg_23_21_inst : DFF_X1 port map( D => N300, CK => clk, Q => n26464, QN
                           => n1973);
   regs_nxt_reg_23_20_inst : DLH_X1 port map( G => n27629, D => n27283, Q => 
                           regs_nxt_23_20_port);
   regs_reg_23_20_inst : DFF_X1 port map( D => N299, CK => clk, Q => n26463, QN
                           => n1969);
   regs_nxt_reg_23_19_inst : DLH_X1 port map( G => n27629, D => n27289, Q => 
                           regs_nxt_23_19_port);
   regs_reg_23_19_inst : DFF_X1 port map( D => N298, CK => clk, Q => n26462, QN
                           => n1965);
   regs_nxt_reg_23_18_inst : DLH_X1 port map( G => n27631, D => n27295, Q => 
                           regs_nxt_23_18_port);
   regs_reg_23_18_inst : DFF_X1 port map( D => N297, CK => clk, Q => n26461, QN
                           => n1961);
   regs_nxt_reg_23_17_inst : DLH_X1 port map( G => n27629, D => n27301, Q => 
                           regs_nxt_23_17_port);
   regs_reg_23_17_inst : DFF_X1 port map( D => N296, CK => clk, Q => n26460, QN
                           => n1957);
   regs_nxt_reg_23_16_inst : DLH_X1 port map( G => n27631, D => n27307, Q => 
                           regs_nxt_23_16_port);
   regs_reg_23_16_inst : DFF_X1 port map( D => N295, CK => clk, Q => n26459, QN
                           => n1953);
   regs_nxt_reg_23_15_inst : DLH_X1 port map( G => n27629, D => n27313, Q => 
                           regs_nxt_23_15_port);
   regs_reg_23_15_inst : DFF_X1 port map( D => N294, CK => clk, Q => n26458, QN
                           => n1949);
   regs_nxt_reg_23_14_inst : DLH_X1 port map( G => n27631, D => n27319, Q => 
                           regs_nxt_23_14_port);
   regs_reg_23_14_inst : DFF_X1 port map( D => N293, CK => clk, Q => n26457, QN
                           => n1945);
   regs_nxt_reg_23_13_inst : DLH_X1 port map( G => n27631, D => n27325, Q => 
                           regs_nxt_23_13_port);
   regs_reg_23_13_inst : DFF_X1 port map( D => N292, CK => clk, Q => n26456, QN
                           => n1941);
   regs_nxt_reg_23_12_inst : DLH_X1 port map( G => n27631, D => n27331, Q => 
                           regs_nxt_23_12_port);
   regs_reg_23_12_inst : DFF_X1 port map( D => N291, CK => clk, Q => n26455, QN
                           => n1937);
   regs_nxt_reg_23_11_inst : DLH_X1 port map( G => n27629, D => n27337, Q => 
                           regs_nxt_23_11_port);
   regs_reg_23_11_inst : DFF_X1 port map( D => N290, CK => clk, Q => n26454, QN
                           => n1933);
   regs_nxt_reg_23_10_inst : DLH_X1 port map( G => n27629, D => n27343, Q => 
                           regs_nxt_23_10_port);
   regs_reg_23_10_inst : DFF_X1 port map( D => N289, CK => clk, Q => n26453, QN
                           => n1929);
   regs_nxt_reg_23_9_inst : DLH_X1 port map( G => n27630, D => n27349, Q => 
                           regs_nxt_23_9_port);
   regs_reg_23_9_inst : DFF_X1 port map( D => N288, CK => clk, Q => n26452, QN 
                           => n1925);
   regs_nxt_reg_23_8_inst : DLH_X1 port map( G => n27630, D => n27357, Q => 
                           regs_nxt_23_8_port);
   regs_reg_23_8_inst : DFF_X1 port map( D => N287, CK => clk, Q => n26451, QN 
                           => n1921);
   regs_nxt_reg_23_7_inst : DLH_X1 port map( G => n27630, D => n27361, Q => 
                           regs_nxt_23_7_port);
   regs_reg_23_7_inst : DFF_X1 port map( D => N286, CK => clk, Q => n26450, QN 
                           => n1917);
   regs_nxt_reg_23_6_inst : DLH_X1 port map( G => n27630, D => n27367, Q => 
                           regs_nxt_23_6_port);
   regs_reg_23_6_inst : DFF_X1 port map( D => N285, CK => clk, Q => n26449, QN 
                           => n1913);
   regs_nxt_reg_23_5_inst : DLH_X1 port map( G => n27630, D => n27277, Q => 
                           regs_nxt_23_5_port);
   regs_reg_23_5_inst : DFF_X1 port map( D => N284, CK => clk, Q => n26448, QN 
                           => n1909);
   regs_nxt_reg_23_4_inst : DLH_X1 port map( G => n27630, D => n27439, Q => 
                           regs_nxt_23_4_port);
   regs_reg_23_4_inst : DFF_X1 port map( D => N283, CK => clk, Q => n26447, QN 
                           => n1905);
   regs_nxt_reg_23_3_inst : DLH_X1 port map( G => n27631, D => n27445, Q => 
                           regs_nxt_23_3_port);
   regs_reg_23_3_inst : DFF_X1 port map( D => N282, CK => clk, Q => n26446, QN 
                           => n1901);
   regs_nxt_reg_23_2_inst : DLH_X1 port map( G => n27630, D => n27451, Q => 
                           regs_nxt_23_2_port);
   regs_reg_23_2_inst : DFF_X1 port map( D => N281, CK => clk, Q => n26445, QN 
                           => n1897);
   regs_nxt_reg_23_1_inst : DLH_X1 port map( G => n27629, D => n27457, Q => 
                           regs_nxt_23_1_port);
   regs_reg_23_1_inst : DFF_X1 port map( D => N280, CK => clk, Q => n26444, QN 
                           => n1893);
   regs_nxt_reg_23_0_inst : DLH_X1 port map( G => n27630, D => n27463, Q => 
                           regs_nxt_23_0_port);
   regs_reg_23_0_inst : DFF_X1 port map( D => N279, CK => clk, Q => n26443, QN 
                           => n1889);
   regs_nxt_reg_24_31_inst : DLH_X1 port map( G => n27637, D => n27373, Q => 
                           regs_nxt_24_31_port);
   regs_reg_24_31_inst : DFF_X1 port map( D => N278, CK => clk, Q => n2221, QN 
                           => n26889);
   regs_nxt_reg_24_30_inst : DLH_X1 port map( G => n27637, D => n27379, Q => 
                           regs_nxt_24_30_port);
   regs_reg_24_30_inst : DFF_X1 port map( D => N277, CK => clk, Q => n2214, QN 
                           => n26887);
   regs_nxt_reg_24_29_inst : DLH_X1 port map( G => n27636, D => n27385, Q => 
                           regs_nxt_24_29_port);
   regs_reg_24_29_inst : DFF_X1 port map( D => N276, CK => clk, Q => n2207, QN 
                           => n26885);
   regs_nxt_reg_24_28_inst : DLH_X1 port map( G => n27636, D => n27391, Q => 
                           regs_nxt_24_28_port);
   regs_reg_24_28_inst : DFF_X1 port map( D => N275, CK => clk, Q => n2200, QN 
                           => n26883);
   regs_nxt_reg_24_27_inst : DLH_X1 port map( G => n27639, D => n27397, Q => 
                           regs_nxt_24_27_port);
   regs_reg_24_27_inst : DFF_X1 port map( D => N274, CK => clk, Q => n2193, QN 
                           => n26881);
   regs_nxt_reg_24_26_inst : DLH_X1 port map( G => n27638, D => n27403, Q => 
                           regs_nxt_24_26_port);
   regs_reg_24_26_inst : DFF_X1 port map( D => N273, CK => clk, Q => n2186, QN 
                           => n26879);
   regs_nxt_reg_24_25_inst : DLH_X1 port map( G => n27639, D => n27409, Q => 
                           regs_nxt_24_25_port);
   regs_reg_24_25_inst : DFF_X1 port map( D => N272, CK => clk, Q => n2179, QN 
                           => n26877);
   regs_nxt_reg_24_24_inst : DLH_X1 port map( G => n27638, D => n27415, Q => 
                           regs_nxt_24_24_port);
   regs_reg_24_24_inst : DFF_X1 port map( D => N271, CK => clk, Q => n2172, QN 
                           => n26875);
   regs_nxt_reg_24_23_inst : DLH_X1 port map( G => n27638, D => n27421, Q => 
                           regs_nxt_24_23_port);
   regs_reg_24_23_inst : DFF_X1 port map( D => N270, CK => clk, Q => n2165, QN 
                           => n26873);
   regs_nxt_reg_24_22_inst : DLH_X1 port map( G => n27638, D => n27427, Q => 
                           regs_nxt_24_22_port);
   regs_reg_24_22_inst : DFF_X1 port map( D => N269, CK => clk, Q => n2158, QN 
                           => n26871);
   regs_nxt_reg_24_21_inst : DLH_X1 port map( G => n27636, D => n27433, Q => 
                           regs_nxt_24_21_port);
   regs_reg_24_21_inst : DFF_X1 port map( D => N268, CK => clk, Q => n2151, QN 
                           => n26869);
   regs_nxt_reg_24_20_inst : DLH_X1 port map( G => n27636, D => n27283, Q => 
                           regs_nxt_24_20_port);
   regs_reg_24_20_inst : DFF_X1 port map( D => N267, CK => clk, Q => n2144, QN 
                           => n26867);
   regs_nxt_reg_24_19_inst : DLH_X1 port map( G => n27636, D => n27289, Q => 
                           regs_nxt_24_19_port);
   regs_reg_24_19_inst : DFF_X1 port map( D => N266, CK => clk, Q => n2137, QN 
                           => n26865);
   regs_nxt_reg_24_18_inst : DLH_X1 port map( G => n27638, D => n27295, Q => 
                           regs_nxt_24_18_port);
   regs_reg_24_18_inst : DFF_X1 port map( D => N265, CK => clk, Q => n2134, QN 
                           => n26864);
   regs_nxt_reg_24_17_inst : DLH_X1 port map( G => n27636, D => n27301, Q => 
                           regs_nxt_24_17_port);
   regs_reg_24_17_inst : DFF_X1 port map( D => N264, CK => clk, Q => n2131, QN 
                           => n26863);
   regs_nxt_reg_24_16_inst : DLH_X1 port map( G => n27638, D => n27307, Q => 
                           regs_nxt_24_16_port);
   regs_reg_24_16_inst : DFF_X1 port map( D => N263, CK => clk, Q => n2128, QN 
                           => n26862);
   regs_nxt_reg_24_15_inst : DLH_X1 port map( G => n27636, D => n27313, Q => 
                           regs_nxt_24_15_port);
   regs_reg_24_15_inst : DFF_X1 port map( D => N262, CK => clk, Q => n2125, QN 
                           => n26861);
   regs_nxt_reg_24_14_inst : DLH_X1 port map( G => n27638, D => n27319, Q => 
                           regs_nxt_24_14_port);
   regs_reg_24_14_inst : DFF_X1 port map( D => N261, CK => clk, Q => n2122, QN 
                           => n26860);
   regs_nxt_reg_24_13_inst : DLH_X1 port map( G => n27638, D => n27325, Q => 
                           regs_nxt_24_13_port);
   regs_reg_24_13_inst : DFF_X1 port map( D => N260, CK => clk, Q => n2119, QN 
                           => n26859);
   regs_nxt_reg_24_12_inst : DLH_X1 port map( G => n27638, D => n27331, Q => 
                           regs_nxt_24_12_port);
   regs_reg_24_12_inst : DFF_X1 port map( D => N259, CK => clk, Q => n2116, QN 
                           => n26858);
   regs_nxt_reg_24_11_inst : DLH_X1 port map( G => n27636, D => n27337, Q => 
                           regs_nxt_24_11_port);
   regs_reg_24_11_inst : DFF_X1 port map( D => N258, CK => clk, Q => n2113, QN 
                           => n26857);
   regs_nxt_reg_24_10_inst : DLH_X1 port map( G => n27636, D => n27343, Q => 
                           regs_nxt_24_10_port);
   regs_reg_24_10_inst : DFF_X1 port map( D => N257, CK => clk, Q => n2110, QN 
                           => n26856);
   regs_nxt_reg_24_9_inst : DLH_X1 port map( G => n27637, D => n27349, Q => 
                           regs_nxt_24_9_port);
   regs_reg_24_9_inst : DFF_X1 port map( D => N256, CK => clk, Q => n2107, QN 
                           => n26855);
   regs_nxt_reg_24_8_inst : DLH_X1 port map( G => n27637, D => n27355, Q => 
                           regs_nxt_24_8_port);
   regs_reg_24_8_inst : DFF_X1 port map( D => N255, CK => clk, Q => n2104, QN 
                           => n26854);
   regs_nxt_reg_24_7_inst : DLH_X1 port map( G => n27637, D => n27361, Q => 
                           regs_nxt_24_7_port);
   regs_reg_24_7_inst : DFF_X1 port map( D => N254, CK => clk, Q => n2101, QN 
                           => n26853);
   regs_nxt_reg_24_6_inst : DLH_X1 port map( G => n27637, D => n27367, Q => 
                           regs_nxt_24_6_port);
   regs_reg_24_6_inst : DFF_X1 port map( D => N253, CK => clk, Q => n2098, QN 
                           => n26852);
   regs_nxt_reg_24_5_inst : DLH_X1 port map( G => n27637, D => n27277, Q => 
                           regs_nxt_24_5_port);
   regs_reg_24_5_inst : DFF_X1 port map( D => N252, CK => clk, Q => n2095, QN 
                           => n26851);
   regs_nxt_reg_24_4_inst : DLH_X1 port map( G => n27637, D => n27439, Q => 
                           regs_nxt_24_4_port);
   regs_reg_24_4_inst : DFF_X1 port map( D => N251, CK => clk, Q => n2092, QN 
                           => n26850);
   regs_nxt_reg_24_3_inst : DLH_X1 port map( G => n27638, D => n27445, Q => 
                           regs_nxt_24_3_port);
   regs_reg_24_3_inst : DFF_X1 port map( D => N250, CK => clk, Q => n2089, QN 
                           => n26849);
   regs_nxt_reg_24_2_inst : DLH_X1 port map( G => n27637, D => n27451, Q => 
                           regs_nxt_24_2_port);
   regs_reg_24_2_inst : DFF_X1 port map( D => N249, CK => clk, Q => n2086, QN 
                           => n26848);
   regs_nxt_reg_24_1_inst : DLH_X1 port map( G => n27636, D => n27457, Q => 
                           regs_nxt_24_1_port);
   regs_reg_24_1_inst : DFF_X1 port map( D => N248, CK => clk, Q => n2083, QN 
                           => n26847);
   regs_nxt_reg_24_0_inst : DLH_X1 port map( G => n27637, D => n27463, Q => 
                           regs_nxt_24_0_port);
   regs_reg_24_0_inst : DFF_X1 port map( D => N247, CK => clk, Q => n2080, QN 
                           => n26846);
   regs_nxt_reg_25_31_inst : DLH_X1 port map( G => n27644, D => n27373, Q => 
                           regs_nxt_25_31_port);
   regs_reg_25_31_inst : DFF_X1 port map( D => N246, CK => clk, Q => n26781, QN
                           => n2612);
   regs_nxt_reg_25_30_inst : DLH_X1 port map( G => n27644, D => n27379, Q => 
                           regs_nxt_25_30_port);
   regs_reg_25_30_inst : DFF_X1 port map( D => N245, CK => clk, Q => n26780, QN
                           => n2608);
   regs_nxt_reg_25_29_inst : DLH_X1 port map( G => n27643, D => n27385, Q => 
                           regs_nxt_25_29_port);
   regs_reg_25_29_inst : DFF_X1 port map( D => N244, CK => clk, Q => n26779, QN
                           => n2604);
   regs_nxt_reg_25_28_inst : DLH_X1 port map( G => n27643, D => n27391, Q => 
                           regs_nxt_25_28_port);
   regs_reg_25_28_inst : DFF_X1 port map( D => N243, CK => clk, Q => n26778, QN
                           => n2600);
   regs_nxt_reg_25_27_inst : DLH_X1 port map( G => n27646, D => n27397, Q => 
                           regs_nxt_25_27_port);
   regs_reg_25_27_inst : DFF_X1 port map( D => N242, CK => clk, Q => n26777, QN
                           => n2596);
   regs_nxt_reg_25_26_inst : DLH_X1 port map( G => n27645, D => n27403, Q => 
                           regs_nxt_25_26_port);
   regs_reg_25_26_inst : DFF_X1 port map( D => N241, CK => clk, Q => n26776, QN
                           => n2592);
   regs_nxt_reg_25_25_inst : DLH_X1 port map( G => n27646, D => n27409, Q => 
                           regs_nxt_25_25_port);
   regs_reg_25_25_inst : DFF_X1 port map( D => N240, CK => clk, Q => n26775, QN
                           => n2588);
   regs_nxt_reg_25_24_inst : DLH_X1 port map( G => n27645, D => n27415, Q => 
                           regs_nxt_25_24_port);
   regs_reg_25_24_inst : DFF_X1 port map( D => N239, CK => clk, Q => n26774, QN
                           => n2584);
   regs_nxt_reg_25_23_inst : DLH_X1 port map( G => n27645, D => n27421, Q => 
                           regs_nxt_25_23_port);
   regs_reg_25_23_inst : DFF_X1 port map( D => N238, CK => clk, Q => n26773, QN
                           => n2580);
   regs_nxt_reg_25_22_inst : DLH_X1 port map( G => n27645, D => n27427, Q => 
                           regs_nxt_25_22_port);
   regs_reg_25_22_inst : DFF_X1 port map( D => N237, CK => clk, Q => n26772, QN
                           => n2576);
   regs_nxt_reg_25_21_inst : DLH_X1 port map( G => n27643, D => n27433, Q => 
                           regs_nxt_25_21_port);
   regs_reg_25_21_inst : DFF_X1 port map( D => N236, CK => clk, Q => n26771, QN
                           => n2572);
   regs_nxt_reg_25_20_inst : DLH_X1 port map( G => n27643, D => n27283, Q => 
                           regs_nxt_25_20_port);
   regs_reg_25_20_inst : DFF_X1 port map( D => N235, CK => clk, Q => n26770, QN
                           => n2568);
   regs_nxt_reg_25_19_inst : DLH_X1 port map( G => n27643, D => n27289, Q => 
                           regs_nxt_25_19_port);
   regs_reg_25_19_inst : DFF_X1 port map( D => N234, CK => clk, Q => n26769, QN
                           => n2564);
   regs_nxt_reg_25_18_inst : DLH_X1 port map( G => n27645, D => n27295, Q => 
                           regs_nxt_25_18_port);
   regs_reg_25_18_inst : DFF_X1 port map( D => N233, CK => clk, Q => n26768, QN
                           => n2560);
   regs_nxt_reg_25_17_inst : DLH_X1 port map( G => n27643, D => n27301, Q => 
                           regs_nxt_25_17_port);
   regs_reg_25_17_inst : DFF_X1 port map( D => N232, CK => clk, Q => n26767, QN
                           => n2556);
   regs_nxt_reg_25_16_inst : DLH_X1 port map( G => n27645, D => n27307, Q => 
                           regs_nxt_25_16_port);
   regs_reg_25_16_inst : DFF_X1 port map( D => N231, CK => clk, Q => n26766, QN
                           => n2552);
   regs_nxt_reg_25_15_inst : DLH_X1 port map( G => n27643, D => n27313, Q => 
                           regs_nxt_25_15_port);
   regs_reg_25_15_inst : DFF_X1 port map( D => N230, CK => clk, Q => n26765, QN
                           => n2548);
   regs_nxt_reg_25_14_inst : DLH_X1 port map( G => n27645, D => n27319, Q => 
                           regs_nxt_25_14_port);
   regs_reg_25_14_inst : DFF_X1 port map( D => N229, CK => clk, Q => n26592, QN
                           => n_1484);
   regs_nxt_reg_25_13_inst : DLH_X1 port map( G => n27645, D => n27325, Q => 
                           regs_nxt_25_13_port);
   regs_reg_25_13_inst : DFF_X1 port map( D => N228, CK => clk, Q => n26591, QN
                           => n_1485);
   regs_nxt_reg_25_12_inst : DLH_X1 port map( G => n27645, D => n27331, Q => 
                           regs_nxt_25_12_port);
   regs_reg_25_12_inst : DFF_X1 port map( D => N227, CK => clk, Q => n26590, QN
                           => n_1486);
   regs_nxt_reg_25_11_inst : DLH_X1 port map( G => n27643, D => n27337, Q => 
                           regs_nxt_25_11_port);
   regs_reg_25_11_inst : DFF_X1 port map( D => N226, CK => clk, Q => n26589, QN
                           => n_1487);
   regs_nxt_reg_25_10_inst : DLH_X1 port map( G => n27643, D => n27343, Q => 
                           regs_nxt_25_10_port);
   regs_reg_25_10_inst : DFF_X1 port map( D => N225, CK => clk, Q => n26595, QN
                           => n_1488);
   regs_nxt_reg_25_9_inst : DLH_X1 port map( G => n27644, D => n27349, Q => 
                           regs_nxt_25_9_port);
   regs_reg_25_9_inst : DFF_X1 port map( D => N224, CK => clk, Q => n26594, QN 
                           => n_1489);
   regs_nxt_reg_25_8_inst : DLH_X1 port map( G => n27644, D => n27355, Q => 
                           regs_nxt_25_8_port);
   regs_reg_25_8_inst : DFF_X1 port map( D => N223, CK => clk, Q => n26593, QN 
                           => n_1490);
   regs_nxt_reg_25_7_inst : DLH_X1 port map( G => n27644, D => n27361, Q => 
                           regs_nxt_25_7_port);
   regs_reg_25_7_inst : DFF_X1 port map( D => N222, CK => clk, Q => n25186, QN 
                           => n_1491);
   regs_nxt_reg_25_6_inst : DLH_X1 port map( G => n27644, D => n27367, Q => 
                           regs_nxt_25_6_port);
   regs_reg_25_6_inst : DFF_X1 port map( D => N221, CK => clk, Q => n25185, QN 
                           => n_1492);
   regs_nxt_reg_25_5_inst : DLH_X1 port map( G => n27644, D => n27277, Q => 
                           regs_nxt_25_5_port);
   regs_reg_25_5_inst : DFF_X1 port map( D => N220, CK => clk, Q => n25184, QN 
                           => n_1493);
   regs_nxt_reg_25_4_inst : DLH_X1 port map( G => n27644, D => n27439, Q => 
                           regs_nxt_25_4_port);
   regs_reg_25_4_inst : DFF_X1 port map( D => N219, CK => clk, Q => n25183, QN 
                           => n_1494);
   regs_nxt_reg_25_3_inst : DLH_X1 port map( G => n27645, D => n27445, Q => 
                           regs_nxt_25_3_port);
   regs_reg_25_3_inst : DFF_X1 port map( D => N218, CK => clk, Q => n25182, QN 
                           => n_1495);
   regs_nxt_reg_25_2_inst : DLH_X1 port map( G => n27644, D => n27451, Q => 
                           regs_nxt_25_2_port);
   regs_reg_25_2_inst : DFF_X1 port map( D => N217, CK => clk, Q => n25181, QN 
                           => n_1496);
   regs_nxt_reg_25_1_inst : DLH_X1 port map( G => n27643, D => n27457, Q => 
                           regs_nxt_25_1_port);
   regs_reg_25_1_inst : DFF_X1 port map( D => N216, CK => clk, Q => n25180, QN 
                           => n_1497);
   regs_nxt_reg_25_0_inst : DLH_X1 port map( G => n27644, D => n27463, Q => 
                           regs_nxt_25_0_port);
   regs_reg_25_0_inst : DFF_X1 port map( D => N215, CK => clk, Q => n25179, QN 
                           => n_1498);
   regs_nxt_reg_26_31_inst : DLH_X1 port map( G => n27651, D => n27373, Q => 
                           regs_nxt_26_31_port);
   regs_reg_26_31_inst : DFF_X1 port map( D => N214, CK => clk, Q => n2485, QN 
                           => n_1499);
   regs_nxt_reg_26_30_inst : DLH_X1 port map( G => n27651, D => n27379, Q => 
                           regs_nxt_26_30_port);
   regs_reg_26_30_inst : DFF_X1 port map( D => N213, CK => clk, Q => n2483, QN 
                           => n_1500);
   regs_nxt_reg_26_29_inst : DLH_X1 port map( G => n27650, D => n27385, Q => 
                           regs_nxt_26_29_port);
   regs_reg_26_29_inst : DFF_X1 port map( D => N212, CK => clk, Q => n2481, QN 
                           => n_1501);
   regs_nxt_reg_26_28_inst : DLH_X1 port map( G => n27650, D => n27391, Q => 
                           regs_nxt_26_28_port);
   regs_reg_26_28_inst : DFF_X1 port map( D => N211, CK => clk, Q => n2479, QN 
                           => n_1502);
   regs_nxt_reg_26_27_inst : DLH_X1 port map( G => n27653, D => n27397, Q => 
                           regs_nxt_26_27_port);
   regs_reg_26_27_inst : DFF_X1 port map( D => N210, CK => clk, Q => n2477, QN 
                           => n_1503);
   regs_nxt_reg_26_26_inst : DLH_X1 port map( G => n27652, D => n27403, Q => 
                           regs_nxt_26_26_port);
   regs_reg_26_26_inst : DFF_X1 port map( D => N209, CK => clk, Q => n2475, QN 
                           => n_1504);
   regs_nxt_reg_26_25_inst : DLH_X1 port map( G => n27653, D => n27409, Q => 
                           regs_nxt_26_25_port);
   regs_reg_26_25_inst : DFF_X1 port map( D => N208, CK => clk, Q => n2473, QN 
                           => n_1505);
   regs_nxt_reg_26_24_inst : DLH_X1 port map( G => n27652, D => n27415, Q => 
                           regs_nxt_26_24_port);
   regs_reg_26_24_inst : DFF_X1 port map( D => N207, CK => clk, Q => n2471, QN 
                           => n_1506);
   regs_nxt_reg_26_23_inst : DLH_X1 port map( G => n27652, D => n27421, Q => 
                           regs_nxt_26_23_port);
   regs_reg_26_23_inst : DFF_X1 port map( D => N206, CK => clk, Q => n2469, QN 
                           => n_1507);
   regs_nxt_reg_26_22_inst : DLH_X1 port map( G => n27652, D => n27427, Q => 
                           regs_nxt_26_22_port);
   regs_reg_26_22_inst : DFF_X1 port map( D => N205, CK => clk, Q => n2467, QN 
                           => n_1508);
   regs_nxt_reg_26_21_inst : DLH_X1 port map( G => n27650, D => n27433, Q => 
                           regs_nxt_26_21_port);
   regs_reg_26_21_inst : DFF_X1 port map( D => N204, CK => clk, Q => n2465, QN 
                           => n_1509);
   regs_nxt_reg_26_20_inst : DLH_X1 port map( G => n27650, D => n27283, Q => 
                           regs_nxt_26_20_port);
   regs_reg_26_20_inst : DFF_X1 port map( D => N203, CK => clk, Q => n2463, QN 
                           => n_1510);
   regs_nxt_reg_26_19_inst : DLH_X1 port map( G => n27650, D => n27289, Q => 
                           regs_nxt_26_19_port);
   regs_reg_26_19_inst : DFF_X1 port map( D => N202, CK => clk, Q => n2461, QN 
                           => n_1511);
   regs_nxt_reg_26_18_inst : DLH_X1 port map( G => n27652, D => n27295, Q => 
                           regs_nxt_26_18_port);
   regs_reg_26_18_inst : DFF_X1 port map( D => N201, CK => clk, Q => n2459, QN 
                           => n_1512);
   regs_nxt_reg_26_17_inst : DLH_X1 port map( G => n27650, D => n27301, Q => 
                           regs_nxt_26_17_port);
   regs_reg_26_17_inst : DFF_X1 port map( D => N200, CK => clk, Q => n2457, QN 
                           => n_1513);
   regs_nxt_reg_26_16_inst : DLH_X1 port map( G => n27652, D => n27307, Q => 
                           regs_nxt_26_16_port);
   regs_reg_26_16_inst : DFF_X1 port map( D => N199, CK => clk, Q => n2455_port
                           , QN => n_1514);
   regs_nxt_reg_26_15_inst : DLH_X1 port map( G => n27650, D => n27313, Q => 
                           regs_nxt_26_15_port);
   regs_reg_26_15_inst : DFF_X1 port map( D => N198, CK => clk, Q => n2453, QN 
                           => n_1515);
   regs_nxt_reg_26_14_inst : DLH_X1 port map( G => n27652, D => n27319, Q => 
                           regs_nxt_26_14_port);
   regs_reg_26_14_inst : DFF_X1 port map( D => N197, CK => clk, Q => n2451, QN 
                           => n_1516);
   regs_nxt_reg_26_13_inst : DLH_X1 port map( G => n27652, D => n27325, Q => 
                           regs_nxt_26_13_port);
   regs_reg_26_13_inst : DFF_X1 port map( D => N196, CK => clk, Q => n2449, QN 
                           => n_1517);
   regs_nxt_reg_26_12_inst : DLH_X1 port map( G => n27652, D => n27331, Q => 
                           regs_nxt_26_12_port);
   regs_reg_26_12_inst : DFF_X1 port map( D => N195, CK => clk, Q => n2447, QN 
                           => n_1518);
   regs_nxt_reg_26_11_inst : DLH_X1 port map( G => n27650, D => n27337, Q => 
                           regs_nxt_26_11_port);
   regs_reg_26_11_inst : DFF_X1 port map( D => N194, CK => clk, Q => n2445, QN 
                           => n_1519);
   regs_nxt_reg_26_10_inst : DLH_X1 port map( G => n27650, D => n27343, Q => 
                           regs_nxt_26_10_port);
   regs_reg_26_10_inst : DFF_X1 port map( D => N193, CK => clk, Q => n2443, QN 
                           => n_1520);
   regs_nxt_reg_26_9_inst : DLH_X1 port map( G => n27651, D => n27349, Q => 
                           regs_nxt_26_9_port);
   regs_reg_26_9_inst : DFF_X1 port map( D => N192, CK => clk, Q => n2441, QN 
                           => n_1521);
   regs_nxt_reg_26_8_inst : DLH_X1 port map( G => n27651, D => n27355, Q => 
                           regs_nxt_26_8_port);
   regs_reg_26_8_inst : DFF_X1 port map( D => N191, CK => clk, Q => n2439, QN 
                           => n_1522);
   regs_nxt_reg_26_7_inst : DLH_X1 port map( G => n27651, D => n27361, Q => 
                           regs_nxt_26_7_port);
   regs_reg_26_7_inst : DFF_X1 port map( D => N190, CK => clk, Q => n2437, QN 
                           => n_1523);
   regs_nxt_reg_26_6_inst : DLH_X1 port map( G => n27651, D => n27367, Q => 
                           regs_nxt_26_6_port);
   regs_reg_26_6_inst : DFF_X1 port map( D => N189, CK => clk, Q => n2435, QN 
                           => n_1524);
   regs_nxt_reg_26_5_inst : DLH_X1 port map( G => n27651, D => n27277, Q => 
                           regs_nxt_26_5_port);
   regs_reg_26_5_inst : DFF_X1 port map( D => N188, CK => clk, Q => n2433, QN 
                           => n_1525);
   regs_nxt_reg_26_4_inst : DLH_X1 port map( G => n27651, D => n27439, Q => 
                           regs_nxt_26_4_port);
   regs_reg_26_4_inst : DFF_X1 port map( D => N187, CK => clk, Q => n2431, QN 
                           => n_1526);
   regs_nxt_reg_26_3_inst : DLH_X1 port map( G => n27652, D => n27445, Q => 
                           regs_nxt_26_3_port);
   regs_reg_26_3_inst : DFF_X1 port map( D => N186, CK => clk, Q => n2429, QN 
                           => n_1527);
   regs_nxt_reg_26_2_inst : DLH_X1 port map( G => n27651, D => n27451, Q => 
                           regs_nxt_26_2_port);
   regs_reg_26_2_inst : DFF_X1 port map( D => N185, CK => clk, Q => n2427, QN 
                           => n_1528);
   regs_nxt_reg_26_1_inst : DLH_X1 port map( G => n27650, D => n27457, Q => 
                           regs_nxt_26_1_port);
   regs_reg_26_1_inst : DFF_X1 port map( D => N184, CK => clk, Q => n2425, QN 
                           => n_1529);
   regs_nxt_reg_26_0_inst : DLH_X1 port map( G => n27651, D => n27463, Q => 
                           regs_nxt_26_0_port);
   regs_reg_26_0_inst : DFF_X1 port map( D => N183, CK => clk, Q => n2423_port,
                           QN => n_1530);
   regs_nxt_reg_27_31_inst : DLH_X1 port map( G => n27658, D => n27373, Q => 
                           regs_nxt_27_31_port);
   regs_reg_27_31_inst : DFF_X1 port map( D => N182, CK => clk, Q => n_1531, QN
                           => n2421);
   regs_nxt_reg_27_30_inst : DLH_X1 port map( G => n27658, D => n27379, Q => 
                           regs_nxt_27_30_port);
   regs_reg_27_30_inst : DFF_X1 port map( D => N181, CK => clk, Q => n_1532, QN
                           => n2419);
   regs_nxt_reg_27_29_inst : DLH_X1 port map( G => n27657, D => n27385, Q => 
                           regs_nxt_27_29_port);
   regs_reg_27_29_inst : DFF_X1 port map( D => N180, CK => clk, Q => n_1533, QN
                           => n2417);
   regs_nxt_reg_27_28_inst : DLH_X1 port map( G => n27657, D => n27391, Q => 
                           regs_nxt_27_28_port);
   regs_reg_27_28_inst : DFF_X1 port map( D => N179, CK => clk, Q => n_1534, QN
                           => n2415);
   regs_nxt_reg_27_27_inst : DLH_X1 port map( G => n27660, D => n27397, Q => 
                           regs_nxt_27_27_port);
   regs_reg_27_27_inst : DFF_X1 port map( D => N178, CK => clk, Q => n_1535, QN
                           => n2413);
   regs_nxt_reg_27_26_inst : DLH_X1 port map( G => n27659, D => n27403, Q => 
                           regs_nxt_27_26_port);
   regs_reg_27_26_inst : DFF_X1 port map( D => N177, CK => clk, Q => n_1536, QN
                           => n2411);
   regs_nxt_reg_27_25_inst : DLH_X1 port map( G => n27660, D => n27409, Q => 
                           regs_nxt_27_25_port);
   regs_reg_27_25_inst : DFF_X1 port map( D => N176, CK => clk, Q => n_1537, QN
                           => n2409);
   regs_nxt_reg_27_24_inst : DLH_X1 port map( G => n27659, D => n27415, Q => 
                           regs_nxt_27_24_port);
   regs_reg_27_24_inst : DFF_X1 port map( D => N175, CK => clk, Q => n_1538, QN
                           => n2407);
   regs_nxt_reg_27_23_inst : DLH_X1 port map( G => n27659, D => n27421, Q => 
                           regs_nxt_27_23_port);
   regs_reg_27_23_inst : DFF_X1 port map( D => N174, CK => clk, Q => n_1539, QN
                           => n2405);
   regs_nxt_reg_27_22_inst : DLH_X1 port map( G => n27659, D => n27427, Q => 
                           regs_nxt_27_22_port);
   regs_reg_27_22_inst : DFF_X1 port map( D => N173, CK => clk, Q => n_1540, QN
                           => n2403);
   regs_nxt_reg_27_21_inst : DLH_X1 port map( G => n27657, D => n27433, Q => 
                           regs_nxt_27_21_port);
   regs_reg_27_21_inst : DFF_X1 port map( D => N172, CK => clk, Q => n_1541, QN
                           => n2401);
   regs_nxt_reg_27_20_inst : DLH_X1 port map( G => n27657, D => n27283, Q => 
                           regs_nxt_27_20_port);
   regs_reg_27_20_inst : DFF_X1 port map( D => N171, CK => clk, Q => n_1542, QN
                           => n2399);
   regs_nxt_reg_27_19_inst : DLH_X1 port map( G => n27657, D => n27289, Q => 
                           regs_nxt_27_19_port);
   regs_reg_27_19_inst : DFF_X1 port map( D => N170, CK => clk, Q => n_1543, QN
                           => n2397);
   regs_nxt_reg_27_18_inst : DLH_X1 port map( G => n27659, D => n27295, Q => 
                           regs_nxt_27_18_port);
   regs_reg_27_18_inst : DFF_X1 port map( D => N169, CK => clk, Q => n_1544, QN
                           => n2395);
   regs_nxt_reg_27_17_inst : DLH_X1 port map( G => n27657, D => n27301, Q => 
                           regs_nxt_27_17_port);
   regs_reg_27_17_inst : DFF_X1 port map( D => N168, CK => clk, Q => n_1545, QN
                           => n2393);
   regs_nxt_reg_27_16_inst : DLH_X1 port map( G => n27659, D => n27307, Q => 
                           regs_nxt_27_16_port);
   regs_reg_27_16_inst : DFF_X1 port map( D => N167, CK => clk, Q => n_1546, QN
                           => n2391_port);
   regs_nxt_reg_27_15_inst : DLH_X1 port map( G => n27657, D => n27313, Q => 
                           regs_nxt_27_15_port);
   regs_reg_27_15_inst : DFF_X1 port map( D => N166, CK => clk, Q => n_1547, QN
                           => n2389);
   regs_nxt_reg_27_14_inst : DLH_X1 port map( G => n27659, D => n27319, Q => 
                           regs_nxt_27_14_port);
   regs_reg_27_14_inst : DFF_X1 port map( D => N165, CK => clk, Q => n_1548, QN
                           => n2387);
   regs_nxt_reg_27_13_inst : DLH_X1 port map( G => n27659, D => n27325, Q => 
                           regs_nxt_27_13_port);
   regs_reg_27_13_inst : DFF_X1 port map( D => N164, CK => clk, Q => n_1549, QN
                           => n2385);
   regs_nxt_reg_27_12_inst : DLH_X1 port map( G => n27659, D => n27331, Q => 
                           regs_nxt_27_12_port);
   regs_reg_27_12_inst : DFF_X1 port map( D => N163, CK => clk, Q => n_1550, QN
                           => n2383);
   regs_nxt_reg_27_11_inst : DLH_X1 port map( G => n27657, D => n27337, Q => 
                           regs_nxt_27_11_port);
   regs_reg_27_11_inst : DFF_X1 port map( D => N162, CK => clk, Q => n_1551, QN
                           => n2381);
   regs_nxt_reg_27_10_inst : DLH_X1 port map( G => n27657, D => n27343, Q => 
                           regs_nxt_27_10_port);
   regs_reg_27_10_inst : DFF_X1 port map( D => N161, CK => clk, Q => n_1552, QN
                           => n2379);
   regs_nxt_reg_27_9_inst : DLH_X1 port map( G => n27658, D => n27349, Q => 
                           regs_nxt_27_9_port);
   regs_reg_27_9_inst : DFF_X1 port map( D => N160, CK => clk, Q => n_1553, QN 
                           => n2377);
   regs_nxt_reg_27_8_inst : DLH_X1 port map( G => n27658, D => n27355, Q => 
                           regs_nxt_27_8_port);
   regs_reg_27_8_inst : DFF_X1 port map( D => N159, CK => clk, Q => n_1554, QN 
                           => n2375);
   regs_nxt_reg_27_7_inst : DLH_X1 port map( G => n27658, D => n27361, Q => 
                           regs_nxt_27_7_port);
   regs_reg_27_7_inst : DFF_X1 port map( D => N158, CK => clk, Q => n_1555, QN 
                           => n2373);
   regs_nxt_reg_27_6_inst : DLH_X1 port map( G => n27658, D => n27367, Q => 
                           regs_nxt_27_6_port);
   regs_reg_27_6_inst : DFF_X1 port map( D => N157, CK => clk, Q => n_1556, QN 
                           => n2371);
   regs_nxt_reg_27_5_inst : DLH_X1 port map( G => n27658, D => n27277, Q => 
                           regs_nxt_27_5_port);
   regs_reg_27_5_inst : DFF_X1 port map( D => N156, CK => clk, Q => n_1557, QN 
                           => n2369);
   regs_nxt_reg_27_4_inst : DLH_X1 port map( G => n27658, D => n27439, Q => 
                           regs_nxt_27_4_port);
   regs_reg_27_4_inst : DFF_X1 port map( D => N155, CK => clk, Q => n_1558, QN 
                           => n2367);
   regs_nxt_reg_27_3_inst : DLH_X1 port map( G => n27659, D => n27445, Q => 
                           regs_nxt_27_3_port);
   regs_reg_27_3_inst : DFF_X1 port map( D => N154, CK => clk, Q => n_1559, QN 
                           => n2365);
   regs_nxt_reg_27_2_inst : DLH_X1 port map( G => n27658, D => n27451, Q => 
                           regs_nxt_27_2_port);
   regs_reg_27_2_inst : DFF_X1 port map( D => N153, CK => clk, Q => n_1560, QN 
                           => n2363);
   regs_nxt_reg_27_1_inst : DLH_X1 port map( G => n27657, D => n27457, Q => 
                           regs_nxt_27_1_port);
   regs_reg_27_1_inst : DFF_X1 port map( D => N152, CK => clk, Q => n_1561, QN 
                           => n2361);
   regs_nxt_reg_27_0_inst : DLH_X1 port map( G => n27658, D => n27463, Q => 
                           regs_nxt_27_0_port);
   regs_reg_27_0_inst : DFF_X1 port map( D => N151, CK => clk, Q => n_1562, QN 
                           => n2359_port);
   regs_nxt_reg_28_31_inst : DLH_X1 port map( G => n27665, D => n27373, Q => 
                           regs_nxt_28_31_port);
   regs_reg_28_31_inst : DFF_X1 port map( D => N150, CK => clk, Q => n_1563, QN
                           => n2422);
   regs_nxt_reg_28_30_inst : DLH_X1 port map( G => n27665, D => n27379, Q => 
                           regs_nxt_28_30_port);
   regs_reg_28_30_inst : DFF_X1 port map( D => N149, CK => clk, Q => n_1564, QN
                           => n2420);
   regs_nxt_reg_28_29_inst : DLH_X1 port map( G => n27664, D => n27385, Q => 
                           regs_nxt_28_29_port);
   regs_reg_28_29_inst : DFF_X1 port map( D => N148, CK => clk, Q => n_1565, QN
                           => n2418);
   regs_nxt_reg_28_28_inst : DLH_X1 port map( G => n27664, D => n27391, Q => 
                           regs_nxt_28_28_port);
   regs_reg_28_28_inst : DFF_X1 port map( D => N147, CK => clk, Q => n_1566, QN
                           => n2416);
   regs_nxt_reg_28_27_inst : DLH_X1 port map( G => n27667, D => n27397, Q => 
                           regs_nxt_28_27_port);
   regs_reg_28_27_inst : DFF_X1 port map( D => N146, CK => clk, Q => n_1567, QN
                           => n2414);
   regs_nxt_reg_28_26_inst : DLH_X1 port map( G => n27666, D => n27403, Q => 
                           regs_nxt_28_26_port);
   regs_reg_28_26_inst : DFF_X1 port map( D => N145, CK => clk, Q => n_1568, QN
                           => n2412);
   regs_nxt_reg_28_25_inst : DLH_X1 port map( G => n27667, D => n27409, Q => 
                           regs_nxt_28_25_port);
   regs_reg_28_25_inst : DFF_X1 port map( D => N144, CK => clk, Q => n_1569, QN
                           => n2410);
   regs_nxt_reg_28_24_inst : DLH_X1 port map( G => n27666, D => n27415, Q => 
                           regs_nxt_28_24_port);
   regs_reg_28_24_inst : DFF_X1 port map( D => N143, CK => clk, Q => n_1570, QN
                           => n2408);
   regs_nxt_reg_28_23_inst : DLH_X1 port map( G => n27666, D => n27421, Q => 
                           regs_nxt_28_23_port);
   regs_reg_28_23_inst : DFF_X1 port map( D => N142, CK => clk, Q => n_1571, QN
                           => n2406);
   regs_nxt_reg_28_22_inst : DLH_X1 port map( G => n27666, D => n27427, Q => 
                           regs_nxt_28_22_port);
   regs_reg_28_22_inst : DFF_X1 port map( D => N141, CK => clk, Q => n_1572, QN
                           => n2404);
   regs_nxt_reg_28_21_inst : DLH_X1 port map( G => n27664, D => n27433, Q => 
                           regs_nxt_28_21_port);
   regs_reg_28_21_inst : DFF_X1 port map( D => N140, CK => clk, Q => n_1573, QN
                           => n2402);
   regs_nxt_reg_28_20_inst : DLH_X1 port map( G => n27664, D => n27283, Q => 
                           regs_nxt_28_20_port);
   regs_reg_28_20_inst : DFF_X1 port map( D => N139, CK => clk, Q => n_1574, QN
                           => n2400);
   regs_nxt_reg_28_19_inst : DLH_X1 port map( G => n27664, D => n27289, Q => 
                           regs_nxt_28_19_port);
   regs_reg_28_19_inst : DFF_X1 port map( D => N138, CK => clk, Q => n_1575, QN
                           => n2398);
   regs_nxt_reg_28_18_inst : DLH_X1 port map( G => n27666, D => n27295, Q => 
                           regs_nxt_28_18_port);
   regs_reg_28_18_inst : DFF_X1 port map( D => N137, CK => clk, Q => n_1576, QN
                           => n2396);
   regs_nxt_reg_28_17_inst : DLH_X1 port map( G => n27664, D => n27301, Q => 
                           regs_nxt_28_17_port);
   regs_reg_28_17_inst : DFF_X1 port map( D => N136, CK => clk, Q => n_1577, QN
                           => n2394);
   regs_nxt_reg_28_16_inst : DLH_X1 port map( G => n27666, D => n27307, Q => 
                           regs_nxt_28_16_port);
   regs_reg_28_16_inst : DFF_X1 port map( D => N135, CK => clk, Q => n_1578, QN
                           => n2392);
   regs_nxt_reg_28_15_inst : DLH_X1 port map( G => n27664, D => n27313, Q => 
                           regs_nxt_28_15_port);
   regs_reg_28_15_inst : DFF_X1 port map( D => N134, CK => clk, Q => n_1579, QN
                           => n2390);
   regs_nxt_reg_28_14_inst : DLH_X1 port map( G => n27666, D => n27319, Q => 
                           regs_nxt_28_14_port);
   regs_reg_28_14_inst : DFF_X1 port map( D => N133, CK => clk, Q => n_1580, QN
                           => n2388);
   regs_nxt_reg_28_13_inst : DLH_X1 port map( G => n27666, D => n27325, Q => 
                           regs_nxt_28_13_port);
   regs_reg_28_13_inst : DFF_X1 port map( D => N132, CK => clk, Q => n_1581, QN
                           => n2386);
   regs_nxt_reg_28_12_inst : DLH_X1 port map( G => n27666, D => n27331, Q => 
                           regs_nxt_28_12_port);
   regs_reg_28_12_inst : DFF_X1 port map( D => N131, CK => clk, Q => n_1582, QN
                           => n2384);
   regs_nxt_reg_28_11_inst : DLH_X1 port map( G => n27664, D => n27337, Q => 
                           regs_nxt_28_11_port);
   regs_reg_28_11_inst : DFF_X1 port map( D => N130, CK => clk, Q => n_1583, QN
                           => n2382);
   regs_nxt_reg_28_10_inst : DLH_X1 port map( G => n27664, D => n27343, Q => 
                           regs_nxt_28_10_port);
   regs_reg_28_10_inst : DFF_X1 port map( D => N129, CK => clk, Q => n_1584, QN
                           => n2380);
   regs_nxt_reg_28_9_inst : DLH_X1 port map( G => n27665, D => n27349, Q => 
                           regs_nxt_28_9_port);
   regs_reg_28_9_inst : DFF_X1 port map( D => N128, CK => clk, Q => n_1585, QN 
                           => n2378);
   regs_nxt_reg_28_8_inst : DLH_X1 port map( G => n27665, D => n27355, Q => 
                           regs_nxt_28_8_port);
   regs_reg_28_8_inst : DFF_X1 port map( D => N127, CK => clk, Q => n_1586, QN 
                           => n2376);
   regs_nxt_reg_28_7_inst : DLH_X1 port map( G => n27665, D => n27361, Q => 
                           regs_nxt_28_7_port);
   regs_reg_28_7_inst : DFF_X1 port map( D => N126, CK => clk, Q => n_1587, QN 
                           => n2374);
   regs_nxt_reg_28_6_inst : DLH_X1 port map( G => n27665, D => n27367, Q => 
                           regs_nxt_28_6_port);
   regs_reg_28_6_inst : DFF_X1 port map( D => N125, CK => clk, Q => n_1588, QN 
                           => n2372);
   regs_nxt_reg_28_5_inst : DLH_X1 port map( G => n27665, D => n27277, Q => 
                           regs_nxt_28_5_port);
   regs_reg_28_5_inst : DFF_X1 port map( D => N124, CK => clk, Q => n_1589, QN 
                           => n2370);
   regs_nxt_reg_28_4_inst : DLH_X1 port map( G => n27665, D => n27439, Q => 
                           regs_nxt_28_4_port);
   regs_reg_28_4_inst : DFF_X1 port map( D => N123, CK => clk, Q => n_1590, QN 
                           => n2368);
   regs_nxt_reg_28_3_inst : DLH_X1 port map( G => n27666, D => n27445, Q => 
                           regs_nxt_28_3_port);
   regs_reg_28_3_inst : DFF_X1 port map( D => N122, CK => clk, Q => n_1591, QN 
                           => n2366);
   regs_nxt_reg_28_2_inst : DLH_X1 port map( G => n27665, D => n27451, Q => 
                           regs_nxt_28_2_port);
   regs_reg_28_2_inst : DFF_X1 port map( D => N121, CK => clk, Q => n_1592, QN 
                           => n2364);
   regs_nxt_reg_28_1_inst : DLH_X1 port map( G => n27664, D => n27457, Q => 
                           regs_nxt_28_1_port);
   regs_reg_28_1_inst : DFF_X1 port map( D => N120, CK => clk, Q => n_1593, QN 
                           => n2362);
   regs_nxt_reg_28_0_inst : DLH_X1 port map( G => n27665, D => n27463, Q => 
                           regs_nxt_28_0_port);
   regs_reg_28_0_inst : DFF_X1 port map( D => N119, CK => clk, Q => n_1594, QN 
                           => n2360);
   regs_nxt_reg_29_31_inst : DLH_X1 port map( G => n27672, D => n27373, Q => 
                           regs_nxt_29_31_port);
   regs_reg_29_31_inst : DFF_X1 port map( D => N118, CK => clk, Q => n2220, QN 
                           => n26573);
   regs_nxt_reg_29_30_inst : DLH_X1 port map( G => n27672, D => n27379, Q => 
                           regs_nxt_29_30_port);
   regs_reg_29_30_inst : DFF_X1 port map( D => N117, CK => clk, Q => n2213, QN 
                           => n26571);
   regs_nxt_reg_29_29_inst : DLH_X1 port map( G => n27671, D => n27385, Q => 
                           regs_nxt_29_29_port);
   regs_reg_29_29_inst : DFF_X1 port map( D => N116, CK => clk, Q => n2206, QN 
                           => n26569);
   regs_nxt_reg_29_28_inst : DLH_X1 port map( G => n27671, D => n27391, Q => 
                           regs_nxt_29_28_port);
   regs_reg_29_28_inst : DFF_X1 port map( D => N115, CK => clk, Q => n2199_port
                           , QN => n26567);
   regs_nxt_reg_29_27_inst : DLH_X1 port map( G => n27674, D => n27397, Q => 
                           regs_nxt_29_27_port);
   regs_reg_29_27_inst : DFF_X1 port map( D => N114, CK => clk, Q => n2192, QN 
                           => n26565);
   regs_nxt_reg_29_26_inst : DLH_X1 port map( G => n27673, D => n27403, Q => 
                           regs_nxt_29_26_port);
   regs_reg_29_26_inst : DFF_X1 port map( D => N113, CK => clk, Q => n2185, QN 
                           => n26563);
   regs_nxt_reg_29_25_inst : DLH_X1 port map( G => n27674, D => n27409, Q => 
                           regs_nxt_29_25_port);
   regs_reg_29_25_inst : DFF_X1 port map( D => N112, CK => clk, Q => n2178, QN 
                           => n26561);
   regs_nxt_reg_29_24_inst : DLH_X1 port map( G => n27673, D => n27415, Q => 
                           regs_nxt_29_24_port);
   regs_reg_29_24_inst : DFF_X1 port map( D => N111, CK => clk, Q => n2171, QN 
                           => n26559);
   regs_nxt_reg_29_23_inst : DLH_X1 port map( G => n27673, D => n27421, Q => 
                           regs_nxt_29_23_port);
   regs_reg_29_23_inst : DFF_X1 port map( D => N110, CK => clk, Q => n2164, QN 
                           => n26557);
   regs_nxt_reg_29_22_inst : DLH_X1 port map( G => n27673, D => n27427, Q => 
                           regs_nxt_29_22_port);
   regs_reg_29_22_inst : DFF_X1 port map( D => N109, CK => clk, Q => n2157, QN 
                           => n26555);
   regs_nxt_reg_29_21_inst : DLH_X1 port map( G => n27671, D => n27433, Q => 
                           regs_nxt_29_21_port);
   regs_reg_29_21_inst : DFF_X1 port map( D => N108, CK => clk, Q => n2150, QN 
                           => n26553);
   regs_nxt_reg_29_20_inst : DLH_X1 port map( G => n27671, D => n27283, Q => 
                           regs_nxt_29_20_port);
   regs_reg_29_20_inst : DFF_X1 port map( D => N107, CK => clk, Q => n2143, QN 
                           => n26551);
   regs_nxt_reg_29_19_inst : DLH_X1 port map( G => n27671, D => n27289, Q => 
                           regs_nxt_29_19_port);
   regs_reg_29_19_inst : DFF_X1 port map( D => N106, CK => clk, Q => n2136, QN 
                           => n26549);
   regs_nxt_reg_29_18_inst : DLH_X1 port map( G => n27673, D => n27295, Q => 
                           regs_nxt_29_18_port);
   regs_reg_29_18_inst : DFF_X1 port map( D => N105, CK => clk, Q => n2133, QN 
                           => n26548);
   regs_nxt_reg_29_17_inst : DLH_X1 port map( G => n27671, D => n27301, Q => 
                           regs_nxt_29_17_port);
   regs_reg_29_17_inst : DFF_X1 port map( D => N104, CK => clk, Q => n2130, QN 
                           => n26547);
   regs_nxt_reg_29_16_inst : DLH_X1 port map( G => n27673, D => n27307, Q => 
                           regs_nxt_29_16_port);
   regs_reg_29_16_inst : DFF_X1 port map( D => N103, CK => clk, Q => n2127, QN 
                           => n26546);
   regs_nxt_reg_29_15_inst : DLH_X1 port map( G => n27671, D => n27313, Q => 
                           regs_nxt_29_15_port);
   regs_reg_29_15_inst : DFF_X1 port map( D => N102, CK => clk, Q => n2124, QN 
                           => n26545);
   regs_nxt_reg_29_14_inst : DLH_X1 port map( G => n27673, D => n27319, Q => 
                           regs_nxt_29_14_port);
   regs_reg_29_14_inst : DFF_X1 port map( D => N101, CK => clk, Q => n2121, QN 
                           => n26544);
   regs_nxt_reg_29_13_inst : DLH_X1 port map( G => n27673, D => n27325, Q => 
                           regs_nxt_29_13_port);
   regs_reg_29_13_inst : DFF_X1 port map( D => N100, CK => clk, Q => n2118, QN 
                           => n26543);
   regs_nxt_reg_29_12_inst : DLH_X1 port map( G => n27673, D => n27331, Q => 
                           regs_nxt_29_12_port);
   regs_reg_29_12_inst : DFF_X1 port map( D => N99, CK => clk, Q => n2115, QN 
                           => n26542);
   regs_nxt_reg_29_11_inst : DLH_X1 port map( G => n27671, D => n27337, Q => 
                           regs_nxt_29_11_port);
   regs_reg_29_11_inst : DFF_X1 port map( D => N98, CK => clk, Q => n2112, QN 
                           => n26541);
   regs_nxt_reg_29_10_inst : DLH_X1 port map( G => n27671, D => n27343, Q => 
                           regs_nxt_29_10_port);
   regs_reg_29_10_inst : DFF_X1 port map( D => N97, CK => clk, Q => n2109, QN 
                           => n26540);
   regs_nxt_reg_29_9_inst : DLH_X1 port map( G => n27672, D => n27349, Q => 
                           regs_nxt_29_9_port);
   regs_reg_29_9_inst : DFF_X1 port map( D => N96, CK => clk, Q => n2106, QN =>
                           n26539);
   regs_nxt_reg_29_8_inst : DLH_X1 port map( G => n27672, D => n27355, Q => 
                           regs_nxt_29_8_port);
   regs_reg_29_8_inst : DFF_X1 port map( D => N95, CK => clk, Q => n2103, QN =>
                           n26538);
   regs_nxt_reg_29_7_inst : DLH_X1 port map( G => n27672, D => n27361, Q => 
                           regs_nxt_29_7_port);
   regs_reg_29_7_inst : DFF_X1 port map( D => N94, CK => clk, Q => n2100, QN =>
                           n26537);
   regs_nxt_reg_29_6_inst : DLH_X1 port map( G => n27672, D => n27367, Q => 
                           regs_nxt_29_6_port);
   regs_reg_29_6_inst : DFF_X1 port map( D => N93, CK => clk, Q => n2097, QN =>
                           n26536);
   regs_nxt_reg_29_5_inst : DLH_X1 port map( G => n27672, D => n27277, Q => 
                           regs_nxt_29_5_port);
   regs_reg_29_5_inst : DFF_X1 port map( D => N92, CK => clk, Q => n2094, QN =>
                           n26535);
   regs_nxt_reg_29_4_inst : DLH_X1 port map( G => n27672, D => n27439, Q => 
                           regs_nxt_29_4_port);
   regs_reg_29_4_inst : DFF_X1 port map( D => N91, CK => clk, Q => n2091, QN =>
                           n26534);
   regs_nxt_reg_29_3_inst : DLH_X1 port map( G => n27673, D => n27445, Q => 
                           regs_nxt_29_3_port);
   regs_reg_29_3_inst : DFF_X1 port map( D => N90, CK => clk, Q => n2088, QN =>
                           n26533);
   regs_nxt_reg_29_2_inst : DLH_X1 port map( G => n27672, D => n27451, Q => 
                           regs_nxt_29_2_port);
   regs_reg_29_2_inst : DFF_X1 port map( D => N89, CK => clk, Q => n2085, QN =>
                           n26532);
   regs_nxt_reg_29_1_inst : DLH_X1 port map( G => n27671, D => n27457, Q => 
                           regs_nxt_29_1_port);
   regs_reg_29_1_inst : DFF_X1 port map( D => N88, CK => clk, Q => n2082, QN =>
                           n26531);
   regs_nxt_reg_29_0_inst : DLH_X1 port map( G => n27672, D => n27463, Q => 
                           regs_nxt_29_0_port);
   regs_reg_29_0_inst : DFF_X1 port map( D => N87, CK => clk, Q => n2079, QN =>
                           n26530);
   regs_nxt_reg_30_31_inst : DLH_X1 port map( G => n27679, D => n27372, Q => 
                           regs_nxt_30_31_port);
   regs_reg_30_31_inst : DFF_X1 port map( D => N86, CK => clk, Q => n2486, QN 
                           => n_1595);
   regs_nxt_reg_30_30_inst : DLH_X1 port map( G => n27679, D => n27378, Q => 
                           regs_nxt_30_30_port);
   regs_reg_30_30_inst : DFF_X1 port map( D => N85, CK => clk, Q => n2484, QN 
                           => n_1596);
   regs_nxt_reg_30_29_inst : DLH_X1 port map( G => n27678, D => n27384, Q => 
                           regs_nxt_30_29_port);
   regs_reg_30_29_inst : DFF_X1 port map( D => N84, CK => clk, Q => n2482, QN 
                           => n_1597);
   regs_nxt_reg_30_28_inst : DLH_X1 port map( G => n27678, D => n27390, Q => 
                           regs_nxt_30_28_port);
   regs_reg_30_28_inst : DFF_X1 port map( D => N83, CK => clk, Q => n2480, QN 
                           => n_1598);
   regs_nxt_reg_30_27_inst : DLH_X1 port map( G => n27681, D => n27396, Q => 
                           regs_nxt_30_27_port);
   regs_reg_30_27_inst : DFF_X1 port map( D => N82, CK => clk, Q => n2478, QN 
                           => n_1599);
   regs_nxt_reg_30_26_inst : DLH_X1 port map( G => n27680, D => n27402, Q => 
                           regs_nxt_30_26_port);
   regs_reg_30_26_inst : DFF_X1 port map( D => N81, CK => clk, Q => n2476, QN 
                           => n_1600);
   regs_nxt_reg_30_25_inst : DLH_X1 port map( G => n27681, D => n27408, Q => 
                           regs_nxt_30_25_port);
   regs_reg_30_25_inst : DFF_X1 port map( D => N80, CK => clk, Q => n2474, QN 
                           => n_1601);
   regs_nxt_reg_30_24_inst : DLH_X1 port map( G => n27680, D => n27414, Q => 
                           regs_nxt_30_24_port);
   regs_reg_30_24_inst : DFF_X1 port map( D => N79, CK => clk, Q => n2472, QN 
                           => n_1602);
   regs_nxt_reg_30_23_inst : DLH_X1 port map( G => n27680, D => n27420, Q => 
                           regs_nxt_30_23_port);
   regs_reg_30_23_inst : DFF_X1 port map( D => N78, CK => clk, Q => n2470, QN 
                           => n_1603);
   regs_nxt_reg_30_22_inst : DLH_X1 port map( G => n27680, D => n27426, Q => 
                           regs_nxt_30_22_port);
   regs_reg_30_22_inst : DFF_X1 port map( D => N77, CK => clk, Q => n2468, QN 
                           => n_1604);
   regs_nxt_reg_30_21_inst : DLH_X1 port map( G => n27678, D => n27432, Q => 
                           regs_nxt_30_21_port);
   regs_reg_30_21_inst : DFF_X1 port map( D => N76, CK => clk, Q => n2466, QN 
                           => n_1605);
   regs_nxt_reg_30_20_inst : DLH_X1 port map( G => n27678, D => n27282, Q => 
                           regs_nxt_30_20_port);
   regs_reg_30_20_inst : DFF_X1 port map( D => N75, CK => clk, Q => n2464, QN 
                           => n_1606);
   regs_nxt_reg_30_19_inst : DLH_X1 port map( G => n27678, D => n27288, Q => 
                           regs_nxt_30_19_port);
   regs_reg_30_19_inst : DFF_X1 port map( D => N74, CK => clk, Q => n2462, QN 
                           => n_1607);
   regs_nxt_reg_30_18_inst : DLH_X1 port map( G => n27680, D => n27294, Q => 
                           regs_nxt_30_18_port);
   regs_reg_30_18_inst : DFF_X1 port map( D => N73, CK => clk, Q => n2460, QN 
                           => n_1608);
   regs_nxt_reg_30_17_inst : DLH_X1 port map( G => n27678, D => n27300, Q => 
                           regs_nxt_30_17_port);
   regs_reg_30_17_inst : DFF_X1 port map( D => N72, CK => clk, Q => n2458, QN 
                           => n_1609);
   regs_nxt_reg_30_16_inst : DLH_X1 port map( G => n27680, D => n27306, Q => 
                           regs_nxt_30_16_port);
   regs_reg_30_16_inst : DFF_X1 port map( D => N71, CK => clk, Q => n2456, QN 
                           => n_1610);
   regs_nxt_reg_30_15_inst : DLH_X1 port map( G => n27678, D => n27312, Q => 
                           regs_nxt_30_15_port);
   regs_reg_30_15_inst : DFF_X1 port map( D => N70, CK => clk, Q => n2454, QN 
                           => n_1611);
   regs_nxt_reg_30_14_inst : DLH_X1 port map( G => n27680, D => n27318, Q => 
                           regs_nxt_30_14_port);
   regs_reg_30_14_inst : DFF_X1 port map( D => N69, CK => clk, Q => n2452, QN 
                           => n_1612);
   regs_nxt_reg_30_13_inst : DLH_X1 port map( G => n27680, D => n27324, Q => 
                           regs_nxt_30_13_port);
   regs_reg_30_13_inst : DFF_X1 port map( D => N68, CK => clk, Q => n2450, QN 
                           => n_1613);
   regs_nxt_reg_30_12_inst : DLH_X1 port map( G => n27680, D => n27330, Q => 
                           regs_nxt_30_12_port);
   regs_reg_30_12_inst : DFF_X1 port map( D => N67, CK => clk, Q => n2448, QN 
                           => n_1614);
   regs_nxt_reg_30_11_inst : DLH_X1 port map( G => n27678, D => n27336, Q => 
                           regs_nxt_30_11_port);
   regs_reg_30_11_inst : DFF_X1 port map( D => N66, CK => clk, Q => n2446, QN 
                           => n_1615);
   regs_nxt_reg_30_10_inst : DLH_X1 port map( G => n27678, D => n27342, Q => 
                           regs_nxt_30_10_port);
   regs_reg_30_10_inst : DFF_X1 port map( D => N65, CK => clk, Q => n2444, QN 
                           => n_1616);
   regs_nxt_reg_30_9_inst : DLH_X1 port map( G => n27679, D => n27348, Q => 
                           regs_nxt_30_9_port);
   regs_reg_30_9_inst : DFF_X1 port map( D => N64, CK => clk, Q => n2442, QN =>
                           n_1617);
   regs_nxt_reg_30_8_inst : DLH_X1 port map( G => n27679, D => n27355, Q => 
                           regs_nxt_30_8_port);
   regs_reg_30_8_inst : DFF_X1 port map( D => N63, CK => clk, Q => n2440, QN =>
                           n_1618);
   regs_nxt_reg_30_7_inst : DLH_X1 port map( G => n27679, D => n27360, Q => 
                           regs_nxt_30_7_port);
   regs_reg_30_7_inst : DFF_X1 port map( D => N62, CK => clk, Q => n2438, QN =>
                           n_1619);
   regs_nxt_reg_30_6_inst : DLH_X1 port map( G => n27679, D => n27366, Q => 
                           regs_nxt_30_6_port);
   regs_reg_30_6_inst : DFF_X1 port map( D => N61, CK => clk, Q => n2436, QN =>
                           n_1620);
   regs_nxt_reg_30_5_inst : DLH_X1 port map( G => n27679, D => n27276, Q => 
                           regs_nxt_30_5_port);
   regs_reg_30_5_inst : DFF_X1 port map( D => N60, CK => clk, Q => n2434, QN =>
                           n_1621);
   regs_nxt_reg_30_4_inst : DLH_X1 port map( G => n27679, D => n27438, Q => 
                           regs_nxt_30_4_port);
   regs_reg_30_4_inst : DFF_X1 port map( D => N59, CK => clk, Q => n2432, QN =>
                           n_1622);
   regs_nxt_reg_30_3_inst : DLH_X1 port map( G => n27680, D => n27444, Q => 
                           regs_nxt_30_3_port);
   regs_reg_30_3_inst : DFF_X1 port map( D => N58, CK => clk, Q => n2430, QN =>
                           n_1623);
   regs_nxt_reg_30_2_inst : DLH_X1 port map( G => n27679, D => n27450, Q => 
                           regs_nxt_30_2_port);
   regs_reg_30_2_inst : DFF_X1 port map( D => N57, CK => clk, Q => n2428, QN =>
                           n_1624);
   regs_nxt_reg_30_1_inst : DLH_X1 port map( G => n27678, D => n27456, Q => 
                           regs_nxt_30_1_port);
   regs_reg_30_1_inst : DFF_X1 port map( D => N56, CK => clk, Q => n2426, QN =>
                           n_1625);
   regs_nxt_reg_30_0_inst : DLH_X1 port map( G => n27679, D => n27462, Q => 
                           regs_nxt_30_0_port);
   regs_reg_30_0_inst : DFF_X1 port map( D => N55, CK => clk, Q => n2424, QN =>
                           n_1626);
   regs_nxt_reg_31_31_inst : DLH_X1 port map( G => n27686, D => n27375, Q => 
                           regs_nxt_31_31_port);
   regs_reg_31_31_inst : DFF_X1 port map( D => N54, CK => clk, Q => n26729, QN 
                           => n2222);
   regs_nxt_reg_31_30_inst : DLH_X1 port map( G => n27686, D => n27381, Q => 
                           regs_nxt_31_30_port);
   regs_reg_31_30_inst : DFF_X1 port map( D => N53, CK => clk, Q => n26728, QN 
                           => n2215);
   regs_nxt_reg_31_29_inst : DLH_X1 port map( G => n27685, D => n27387, Q => 
                           regs_nxt_31_29_port);
   regs_reg_31_29_inst : DFF_X1 port map( D => N52, CK => clk, Q => n26727, QN 
                           => n2208);
   regs_nxt_reg_31_28_inst : DLH_X1 port map( G => n27685, D => n27393, Q => 
                           regs_nxt_31_28_port);
   regs_reg_31_28_inst : DFF_X1 port map( D => N51, CK => clk, Q => n26726, QN 
                           => n2201);
   regs_nxt_reg_31_27_inst : DLH_X1 port map( G => n27688, D => n27399, Q => 
                           regs_nxt_31_27_port);
   regs_reg_31_27_inst : DFF_X1 port map( D => N50, CK => clk, Q => n26725, QN 
                           => n2194);
   regs_nxt_reg_31_26_inst : DLH_X1 port map( G => n27687, D => n27405, Q => 
                           regs_nxt_31_26_port);
   regs_reg_31_26_inst : DFF_X1 port map( D => N49, CK => clk, Q => n26724, QN 
                           => n2187);
   regs_nxt_reg_31_25_inst : DLH_X1 port map( G => n27688, D => n27411, Q => 
                           regs_nxt_31_25_port);
   regs_reg_31_25_inst : DFF_X1 port map( D => N48, CK => clk, Q => n26723, QN 
                           => n2180);
   regs_nxt_reg_31_24_inst : DLH_X1 port map( G => n27687, D => n27417, Q => 
                           regs_nxt_31_24_port);
   regs_reg_31_24_inst : DFF_X1 port map( D => N47, CK => clk, Q => n26722, QN 
                           => n2173);
   regs_nxt_reg_31_23_inst : DLH_X1 port map( G => n27687, D => n27423, Q => 
                           regs_nxt_31_23_port);
   regs_reg_31_23_inst : DFF_X1 port map( D => N46, CK => clk, Q => n26721, QN 
                           => n2166_port);
   regs_nxt_reg_31_22_inst : DLH_X1 port map( G => n27687, D => n27429, Q => 
                           regs_nxt_31_22_port);
   regs_reg_31_22_inst : DFF_X1 port map( D => N45, CK => clk, Q => n26720, QN 
                           => n2159);
   regs_nxt_reg_31_21_inst : DLH_X1 port map( G => n27685, D => n27435, Q => 
                           regs_nxt_31_21_port);
   regs_reg_31_21_inst : DFF_X1 port map( D => N44, CK => clk, Q => n26719, QN 
                           => n2152);
   regs_nxt_reg_31_20_inst : DLH_X1 port map( G => n27685, D => n27285, Q => 
                           regs_nxt_31_20_port);
   regs_reg_31_20_inst : DFF_X1 port map( D => N43, CK => clk, Q => n26718, QN 
                           => n2145);
   regs_nxt_reg_31_19_inst : DLH_X1 port map( G => n27685, D => n27291, Q => 
                           regs_nxt_31_19_port);
   regs_reg_31_19_inst : DFF_X1 port map( D => N42, CK => clk, Q => n26717, QN 
                           => n2138);
   regs_nxt_reg_31_18_inst : DLH_X1 port map( G => n27687, D => n27297, Q => 
                           regs_nxt_31_18_port);
   regs_reg_31_18_inst : DFF_X1 port map( D => N41, CK => clk, Q => n26716, QN 
                           => n2135);
   regs_nxt_reg_31_17_inst : DLH_X1 port map( G => n27685, D => n27303, Q => 
                           regs_nxt_31_17_port);
   regs_reg_31_17_inst : DFF_X1 port map( D => N40, CK => clk, Q => n26715, QN 
                           => n2132);
   regs_nxt_reg_31_16_inst : DLH_X1 port map( G => n27687, D => n27309, Q => 
                           regs_nxt_31_16_port);
   regs_reg_31_16_inst : DFF_X1 port map( D => N39, CK => clk, Q => n26714, QN 
                           => n2129);
   regs_nxt_reg_31_15_inst : DLH_X1 port map( G => n27685, D => n27315, Q => 
                           regs_nxt_31_15_port);
   regs_reg_31_15_inst : DFF_X1 port map( D => N38, CK => clk, Q => n26713, QN 
                           => n2126);
   regs_nxt_reg_31_14_inst : DLH_X1 port map( G => n27687, D => n27321, Q => 
                           regs_nxt_31_14_port);
   regs_reg_31_14_inst : DFF_X1 port map( D => N37, CK => clk, Q => n26712, QN 
                           => n2123);
   regs_nxt_reg_31_13_inst : DLH_X1 port map( G => n27687, D => n27327, Q => 
                           regs_nxt_31_13_port);
   regs_reg_31_13_inst : DFF_X1 port map( D => N36, CK => clk, Q => n26711, QN 
                           => n2120);
   regs_nxt_reg_31_12_inst : DLH_X1 port map( G => n27687, D => n27333, Q => 
                           regs_nxt_31_12_port);
   regs_reg_31_12_inst : DFF_X1 port map( D => N35, CK => clk, Q => n26710, QN 
                           => n2117);
   regs_nxt_reg_31_11_inst : DLH_X1 port map( G => n27685, D => n27339, Q => 
                           regs_nxt_31_11_port);
   regs_reg_31_11_inst : DFF_X1 port map( D => N34, CK => clk, Q => n26709, QN 
                           => n2114);
   regs_nxt_reg_31_10_inst : DLH_X1 port map( G => n27685, D => n27345, Q => 
                           regs_nxt_31_10_port);
   regs_reg_31_10_inst : DFF_X1 port map( D => N33, CK => clk, Q => n26708, QN 
                           => n2111);
   regs_nxt_reg_31_9_inst : DLH_X1 port map( G => n27686, D => n27351, Q => 
                           regs_nxt_31_9_port);
   regs_reg_31_9_inst : DFF_X1 port map( D => N32, CK => clk, Q => n26707, QN 
                           => n2108);
   regs_nxt_reg_31_8_inst : DLH_X1 port map( G => n27686, D => n27355, Q => 
                           regs_nxt_31_8_port);
   regs_reg_31_8_inst : DFF_X1 port map( D => N31, CK => clk, Q => n26706, QN 
                           => n2105);
   regs_nxt_reg_31_7_inst : DLH_X1 port map( G => n27686, D => n27363, Q => 
                           regs_nxt_31_7_port);
   regs_reg_31_7_inst : DFF_X1 port map( D => N30, CK => clk, Q => n26705, QN 
                           => n2102);
   regs_nxt_reg_31_6_inst : DLH_X1 port map( G => n27686, D => n27369, Q => 
                           regs_nxt_31_6_port);
   regs_reg_31_6_inst : DFF_X1 port map( D => N29, CK => clk, Q => n26704, QN 
                           => n2099);
   regs_nxt_reg_31_5_inst : DLH_X1 port map( G => n27686, D => n27279, Q => 
                           regs_nxt_31_5_port);
   regs_reg_31_5_inst : DFF_X1 port map( D => N28, CK => clk, Q => n26703, QN 
                           => n2096);
   regs_nxt_reg_31_4_inst : DLH_X1 port map( G => n27686, D => n27441, Q => 
                           regs_nxt_31_4_port);
   regs_reg_31_4_inst : DFF_X1 port map( D => N27, CK => clk, Q => n26702, QN 
                           => n2093);
   regs_nxt_reg_31_3_inst : DLH_X1 port map( G => n27687, D => n27447, Q => 
                           regs_nxt_31_3_port);
   regs_reg_31_3_inst : DFF_X1 port map( D => N26, CK => clk, Q => n26701, QN 
                           => n2090);
   regs_nxt_reg_31_2_inst : DLH_X1 port map( G => n27686, D => n27453, Q => 
                           regs_nxt_31_2_port);
   regs_reg_31_2_inst : DFF_X1 port map( D => N25, CK => clk, Q => n26700, QN 
                           => n2087);
   regs_nxt_reg_31_1_inst : DLH_X1 port map( G => n27685, D => n27459, Q => 
                           regs_nxt_31_1_port);
   regs_reg_31_1_inst : DFF_X1 port map( D => N24, CK => clk, Q => n26699, QN 
                           => n2084);
   regs_nxt_reg_31_0_inst : DLH_X1 port map( G => n27686, D => n27465, Q => 
                           regs_nxt_31_0_port);
   regs_reg_31_0_inst : DFF_X1 port map( D => N23, CK => clk, Q => n26698, QN 
                           => n2081);
   U3029 : NAND3_X1 port map( A1 => n27699, A2 => n27700, A3 => wr_en, ZN => 
                           n1875);
   U3030 : NAND3_X1 port map( A1 => wr_en, A2 => n27700, A3 => add_wr(3), ZN =>
                           n1884);
   U3031 : NAND3_X1 port map( A1 => wr_en, A2 => n27699, A3 => add_wr(4), ZN =>
                           n1885);
   U3032 : NAND3_X1 port map( A1 => n27697, A2 => n27698, A3 => n27696, ZN => 
                           n1876);
   U3033 : NAND3_X1 port map( A1 => n27697, A2 => n27698, A3 => add_wr(0), ZN 
                           => n1877);
   U3034 : NAND3_X1 port map( A1 => n27696, A2 => n27698, A3 => add_wr(1), ZN 
                           => n1878);
   U3035 : NAND3_X1 port map( A1 => add_wr(0), A2 => n27698, A3 => add_wr(1), 
                           ZN => n1879);
   U3036 : NAND3_X1 port map( A1 => n27696, A2 => n27697, A3 => add_wr(2), ZN 
                           => n1880);
   U3037 : NAND3_X1 port map( A1 => add_wr(0), A2 => n27697, A3 => add_wr(2), 
                           ZN => n1881);
   U3038 : NAND3_X1 port map( A1 => add_wr(1), A2 => n27696, A3 => add_wr(2), 
                           ZN => n1882);
   U3039 : NAND3_X1 port map( A1 => add_wr(3), A2 => wr_en, A3 => add_wr(4), ZN
                           => n1886);
   U3040 : NAND3_X1 port map( A1 => add_wr(1), A2 => add_wr(0), A3 => add_wr(2)
                           , ZN => n1883);
   U3 : NOR2_X1 port map( A1 => n27714, A2 => add_rd2(4), ZN => n1251);
   U4 : NOR2_X1 port map( A1 => add_rd2(3), A2 => add_rd2(4), ZN => n1250);
   U5 : AND2_X1 port map( A1 => datain(6), A2 => n26996, ZN => n26664);
   U6 : AND2_X1 port map( A1 => datain(7), A2 => n26996, ZN => n26665);
   U7 : AND2_X1 port map( A1 => datain(8), A2 => n26996, ZN => n26666);
   U8 : AND2_X1 port map( A1 => datain(9), A2 => n26996, ZN => n26667);
   U9 : AND2_X1 port map( A1 => datain(10), A2 => n26996, ZN => n26668);
   U10 : AND2_X1 port map( A1 => datain(11), A2 => n26996, ZN => n26669);
   U11 : AND2_X1 port map( A1 => datain(12), A2 => n26996, ZN => n26670);
   U12 : AND2_X1 port map( A1 => datain(13), A2 => n26996, ZN => n26671);
   U13 : AND2_X1 port map( A1 => datain(14), A2 => n26996, ZN => n26672);
   U14 : AND2_X1 port map( A1 => datain(15), A2 => n26996, ZN => n26673);
   U15 : AND2_X1 port map( A1 => datain(16), A2 => n26996, ZN => n26674);
   U16 : AND2_X1 port map( A1 => datain(17), A2 => n26996, ZN => n26675);
   U17 : AND2_X1 port map( A1 => datain(18), A2 => n26996, ZN => n26676);
   U18 : AND2_X1 port map( A1 => datain(19), A2 => n26996, ZN => n26677);
   U19 : AND2_X1 port map( A1 => datain(20), A2 => n26996, ZN => n26678);
   U20 : AND2_X1 port map( A1 => datain(31), A2 => n26996, ZN => n26679);
   U21 : AND2_X1 port map( A1 => datain(0), A2 => n26995, ZN => n26680);
   U22 : AND2_X1 port map( A1 => datain(1), A2 => n26995, ZN => n26681);
   U23 : AND2_X1 port map( A1 => datain(2), A2 => n26995, ZN => n26682);
   U24 : AND2_X1 port map( A1 => datain(3), A2 => n26995, ZN => n26683);
   U25 : AND2_X1 port map( A1 => datain(4), A2 => n26995, ZN => n26684);
   U26 : AND2_X1 port map( A1 => datain(21), A2 => n26995, ZN => n26685);
   U27 : AND2_X1 port map( A1 => datain(22), A2 => n26995, ZN => n26686);
   U28 : AND2_X1 port map( A1 => datain(23), A2 => n26995, ZN => n26687);
   U29 : AND2_X1 port map( A1 => datain(24), A2 => n26995, ZN => n26688);
   U30 : AND2_X1 port map( A1 => datain(25), A2 => n26995, ZN => n26689);
   U31 : AND2_X1 port map( A1 => datain(26), A2 => n26995, ZN => n26690);
   U32 : AND2_X1 port map( A1 => datain(27), A2 => n26995, ZN => n26691);
   U33 : AND2_X1 port map( A1 => datain(28), A2 => n26995, ZN => n26692);
   U34 : AND2_X1 port map( A1 => datain(29), A2 => n26995, ZN => n26693);
   U35 : AND2_X1 port map( A1 => datain(30), A2 => n26995, ZN => n26694);
   U36 : AND2_X1 port map( A1 => datain(5), A2 => n27004, ZN => n26695);
   U37 : BUF_X1 port map( A => n26963, Z => n27191);
   U38 : BUF_X1 port map( A => n26962, Z => n27194);
   U39 : BUF_X1 port map( A => n1293, Z => n27098);
   U40 : BUF_X1 port map( A => n27691, Z => n27689);
   U41 : BUF_X1 port map( A => n27684, Z => n27682);
   U42 : BUF_X1 port map( A => n27677, Z => n27675);
   U43 : BUF_X1 port map( A => n27670, Z => n27668);
   U44 : BUF_X1 port map( A => n27663, Z => n27661);
   U45 : BUF_X1 port map( A => n27656, Z => n27654);
   U46 : BUF_X1 port map( A => n27649, Z => n27647);
   U47 : BUF_X1 port map( A => n27642, Z => n27640);
   U48 : BUF_X1 port map( A => n27635, Z => n27633);
   U49 : BUF_X1 port map( A => n27628, Z => n27626);
   U50 : BUF_X1 port map( A => n27621, Z => n27619);
   U51 : BUF_X1 port map( A => n27614, Z => n27612);
   U52 : BUF_X1 port map( A => n27607, Z => n27605);
   U53 : BUF_X1 port map( A => n27600, Z => n27598);
   U54 : BUF_X1 port map( A => n27593, Z => n27591);
   U55 : BUF_X1 port map( A => n27586, Z => n27584);
   U56 : BUF_X1 port map( A => n27579, Z => n27577);
   U57 : BUF_X1 port map( A => n27572, Z => n27570);
   U58 : BUF_X1 port map( A => n27565, Z => n27563);
   U59 : BUF_X1 port map( A => n27558, Z => n27556);
   U60 : BUF_X1 port map( A => n27551, Z => n27549);
   U61 : BUF_X1 port map( A => n27544, Z => n27542);
   U62 : BUF_X1 port map( A => n27537, Z => n27535);
   U63 : BUF_X1 port map( A => n27530, Z => n27528);
   U64 : BUF_X1 port map( A => n27523, Z => n27521);
   U65 : BUF_X1 port map( A => n27516, Z => n27514);
   U66 : BUF_X1 port map( A => n27509, Z => n27507);
   U67 : BUF_X1 port map( A => n27502, Z => n27500);
   U68 : BUF_X1 port map( A => n27495, Z => n27493);
   U69 : BUF_X1 port map( A => n27488, Z => n27486);
   U70 : BUF_X1 port map( A => n27481, Z => n27479);
   U71 : BUF_X1 port map( A => n27474, Z => n27472);
   U72 : BUF_X1 port map( A => n27720, Z => n26970);
   U73 : BUF_X1 port map( A => n1280, Z => n27126);
   U74 : BUF_X1 port map( A => n1288, Z => n27114);
   U75 : BUF_X1 port map( A => n1289, Z => n27110);
   U76 : BUF_X1 port map( A => n1294, Z => n27094);
   U77 : BUF_X1 port map( A => n1298, Z => n27082);
   U78 : BUF_X1 port map( A => n1299, Z => n27078);
   U79 : BUF_X1 port map( A => n1303, Z => n27066);
   U80 : BUF_X1 port map( A => n1304, Z => n27062);
   U81 : BUF_X1 port map( A => n647_port, Z => n27252);
   U82 : BUF_X1 port map( A => n655_port, Z => n27236);
   U83 : BUF_X1 port map( A => n654_port, Z => n27240);
   U84 : BUF_X1 port map( A => n1262, Z => n27182);
   U85 : BUF_X1 port map( A => n1261, Z => n27186);
   U86 : BUF_X1 port map( A => n1267, Z => n27166);
   U87 : BUF_X1 port map( A => n1266, Z => n27170);
   U88 : BUF_X1 port map( A => n1272, Z => n27150);
   U89 : BUF_X1 port map( A => n1271, Z => n27154);
   U90 : BUF_X1 port map( A => n1277, Z => n27134);
   U91 : BUF_X1 port map( A => n1276, Z => n27138);
   U92 : BUF_X1 port map( A => n26680, Z => n27466);
   U93 : BUF_X1 port map( A => n26681, Z => n27460);
   U94 : BUF_X1 port map( A => n26682, Z => n27454);
   U95 : BUF_X1 port map( A => n26683, Z => n27448);
   U96 : BUF_X1 port map( A => n26684, Z => n27442);
   U97 : BUF_X1 port map( A => n26695, Z => n27280);
   U98 : BUF_X1 port map( A => n26664, Z => n27370);
   U99 : BUF_X1 port map( A => n26665, Z => n27364);
   U100 : BUF_X1 port map( A => n26666, Z => n27358);
   U101 : BUF_X1 port map( A => n26667, Z => n27352);
   U102 : BUF_X1 port map( A => n26668, Z => n27346);
   U103 : BUF_X1 port map( A => n26669, Z => n27340);
   U104 : BUF_X1 port map( A => n26670, Z => n27334);
   U105 : BUF_X1 port map( A => n26671, Z => n27328);
   U106 : BUF_X1 port map( A => n26672, Z => n27322);
   U107 : BUF_X1 port map( A => n26673, Z => n27316);
   U108 : BUF_X1 port map( A => n26674, Z => n27310);
   U109 : BUF_X1 port map( A => n26675, Z => n27304);
   U110 : BUF_X1 port map( A => n26676, Z => n27298);
   U111 : BUF_X1 port map( A => n26677, Z => n27292);
   U112 : BUF_X1 port map( A => n26678, Z => n27286);
   U113 : BUF_X1 port map( A => n26685, Z => n27436);
   U114 : BUF_X1 port map( A => n26686, Z => n27430);
   U115 : BUF_X1 port map( A => n26687, Z => n27424);
   U116 : BUF_X1 port map( A => n26688, Z => n27418);
   U117 : BUF_X1 port map( A => n26689, Z => n27412);
   U118 : BUF_X1 port map( A => n26690, Z => n27406);
   U119 : BUF_X1 port map( A => n26691, Z => n27400);
   U120 : BUF_X1 port map( A => n26692, Z => n27394);
   U121 : BUF_X1 port map( A => n26693, Z => n27388);
   U122 : BUF_X1 port map( A => n26694, Z => n27382);
   U123 : BUF_X1 port map( A => n26679, Z => n27376);
   U124 : BUF_X1 port map( A => n644_port, Z => n27264);
   U125 : BUF_X1 port map( A => n657_port, Z => n27232);
   U126 : BUF_X1 port map( A => n658_port, Z => n27228);
   U127 : BUF_X1 port map( A => n1264, Z => n27178);
   U128 : BUF_X1 port map( A => n1265, Z => n27174);
   U129 : BUF_X1 port map( A => n1269, Z => n27162);
   U130 : BUF_X1 port map( A => n1270, Z => n27158);
   U131 : BUF_X1 port map( A => n1274, Z => n27146);
   U132 : BUF_X1 port map( A => n1275, Z => n27142);
   U133 : BUF_X1 port map( A => n1279, Z => n27130);
   U134 : BUF_X1 port map( A => n642_port, Z => n27268);
   U135 : BUF_X1 port map( A => n641_port, Z => n27272);
   U136 : BUF_X1 port map( A => n646_port, Z => n27256);
   U137 : BUF_X1 port map( A => n664_port, Z => n27220);
   U138 : BUF_X1 port map( A => n663_port, Z => n27224);
   U139 : BUF_X1 port map( A => n669_port, Z => n27204);
   U140 : BUF_X1 port map( A => n668_port, Z => n27208);
   U141 : BUF_X1 port map( A => n1286, Z => n27118);
   U142 : BUF_X1 port map( A => n1285, Z => n27122);
   U143 : BUF_X1 port map( A => n1291, Z => n27102);
   U144 : BUF_X1 port map( A => n1290, Z => n27106);
   U145 : BUF_X1 port map( A => n1296, Z => n27086);
   U146 : BUF_X1 port map( A => n1295, Z => n27090);
   U147 : BUF_X1 port map( A => n1301, Z => n27070);
   U148 : BUF_X1 port map( A => n1300, Z => n27074);
   U149 : BUF_X1 port map( A => n645_port, Z => n27260);
   U150 : BUF_X1 port map( A => n649_port, Z => n27248);
   U151 : BUF_X1 port map( A => n650_port, Z => n27244);
   U152 : BUF_X1 port map( A => n666_port, Z => n27216);
   U153 : BUF_X1 port map( A => n667_port, Z => n27212);
   U154 : BUF_X1 port map( A => n671_port, Z => n27200);
   U155 : BUF_X1 port map( A => n672_port, Z => n27196);
   U156 : BUF_X1 port map( A => n27046, Z => n26995);
   U157 : BUF_X1 port map( A => n27039, Z => n27016);
   U158 : BUF_X1 port map( A => n27039, Z => n27017);
   U159 : BUF_X1 port map( A => n27043, Z => n27005);
   U160 : BUF_X1 port map( A => n27043, Z => n27006);
   U161 : BUF_X1 port map( A => n27042, Z => n27007);
   U162 : BUF_X1 port map( A => n27042, Z => n27008);
   U163 : BUF_X1 port map( A => n27042, Z => n27009);
   U164 : BUF_X1 port map( A => n27041, Z => n27010);
   U165 : BUF_X1 port map( A => n27036, Z => n27027);
   U166 : BUF_X1 port map( A => n27035, Z => n27028);
   U167 : BUF_X1 port map( A => n27035, Z => n27029);
   U168 : BUF_X1 port map( A => n27035, Z => n27030);
   U169 : BUF_X1 port map( A => n27034, Z => n27031);
   U170 : BUF_X1 port map( A => n27034, Z => n27032);
   U171 : BUF_X1 port map( A => n27038, Z => n27019);
   U172 : BUF_X1 port map( A => n27038, Z => n27020);
   U173 : BUF_X1 port map( A => n27038, Z => n27021);
   U174 : BUF_X1 port map( A => n27037, Z => n27022);
   U175 : BUF_X1 port map( A => n27037, Z => n27023);
   U176 : BUF_X1 port map( A => n27037, Z => n27024);
   U177 : BUF_X1 port map( A => n27036, Z => n27025);
   U178 : BUF_X1 port map( A => n27036, Z => n27026);
   U179 : BUF_X1 port map( A => n27051, Z => n26982);
   U180 : BUF_X1 port map( A => n27050, Z => n26983);
   U181 : BUF_X1 port map( A => n27050, Z => n26984);
   U182 : BUF_X1 port map( A => n27050, Z => n26985);
   U183 : BUF_X1 port map( A => n27049, Z => n26986);
   U184 : BUF_X1 port map( A => n27049, Z => n26987);
   U185 : BUF_X1 port map( A => n27049, Z => n26988);
   U186 : BUF_X1 port map( A => n27053, Z => n26975);
   U187 : BUF_X1 port map( A => n27053, Z => n26976);
   U188 : BUF_X1 port map( A => n27052, Z => n26977);
   U189 : BUF_X1 port map( A => n27052, Z => n26978);
   U190 : BUF_X1 port map( A => n27052, Z => n26979);
   U191 : BUF_X1 port map( A => n27051, Z => n26980);
   U192 : BUF_X1 port map( A => n27051, Z => n26981);
   U193 : BUF_X1 port map( A => n27046, Z => n26996);
   U194 : BUF_X1 port map( A => n27046, Z => n26997);
   U195 : BUF_X1 port map( A => n27045, Z => n26998);
   U196 : BUF_X1 port map( A => n27045, Z => n26999);
   U197 : BUF_X1 port map( A => n27045, Z => n27000);
   U198 : BUF_X1 port map( A => n27044, Z => n27001);
   U199 : BUF_X1 port map( A => n27044, Z => n27002);
   U200 : BUF_X1 port map( A => n27044, Z => n27003);
   U201 : BUF_X1 port map( A => n27043, Z => n27004);
   U202 : BUF_X1 port map( A => n27048, Z => n26989);
   U203 : BUF_X1 port map( A => n27048, Z => n26990);
   U204 : BUF_X1 port map( A => n27048, Z => n26991);
   U205 : BUF_X1 port map( A => n27047, Z => n26992);
   U206 : BUF_X1 port map( A => n27047, Z => n26993);
   U207 : BUF_X1 port map( A => n27047, Z => n26994);
   U208 : BUF_X1 port map( A => n27039, Z => n27018);
   U209 : BUF_X1 port map( A => n27040, Z => n27015);
   U210 : BUF_X1 port map( A => n27041, Z => n27011);
   U211 : BUF_X1 port map( A => n27041, Z => n27012);
   U212 : BUF_X1 port map( A => n27040, Z => n27013);
   U213 : BUF_X1 port map( A => n27040, Z => n27014);
   U214 : BUF_X1 port map( A => n27053, Z => n26974);
   U215 : BUF_X1 port map( A => n27054, Z => n26973);
   U216 : BUF_X1 port map( A => n27054, Z => n26972);
   U217 : BUF_X1 port map( A => n27034, Z => n27033);
   U218 : BUF_X1 port map( A => n27057, Z => n27046);
   U219 : BUF_X1 port map( A => n27059, Z => n27042);
   U220 : BUF_X1 port map( A => n27061, Z => n27035);
   U221 : BUF_X1 port map( A => n27061, Z => n27034);
   U222 : BUF_X1 port map( A => n27060, Z => n27038);
   U223 : BUF_X1 port map( A => n27060, Z => n27037);
   U224 : BUF_X1 port map( A => n27061, Z => n27036);
   U225 : BUF_X1 port map( A => n27056, Z => n27050);
   U226 : BUF_X1 port map( A => n27056, Z => n27049);
   U227 : BUF_X1 port map( A => n27055, Z => n27053);
   U228 : BUF_X1 port map( A => n27055, Z => n27052);
   U229 : BUF_X1 port map( A => n27056, Z => n27051);
   U230 : BUF_X1 port map( A => n27058, Z => n27045);
   U231 : BUF_X1 port map( A => n27058, Z => n27044);
   U232 : BUF_X1 port map( A => n27058, Z => n27043);
   U233 : BUF_X1 port map( A => n27057, Z => n27048);
   U234 : BUF_X1 port map( A => n27057, Z => n27047);
   U235 : BUF_X1 port map( A => n27060, Z => n27039);
   U236 : BUF_X1 port map( A => n27059, Z => n27041);
   U237 : BUF_X1 port map( A => n27059, Z => n27040);
   U238 : BUF_X1 port map( A => n27055, Z => n27054);
   U239 : BUF_X1 port map( A => n27098, Z => n27099);
   U240 : BUF_X1 port map( A => n27098, Z => n27100);
   U241 : BUF_X1 port map( A => n27098, Z => n27101);
   U242 : INV_X1 port map( A => n27191, ZN => n27190);
   U243 : INV_X1 port map( A => n27194, ZN => n27193);
   U244 : BUF_X1 port map( A => n27689, Z => n27687);
   U245 : BUF_X1 port map( A => n27689, Z => n27686);
   U246 : BUF_X1 port map( A => n27682, Z => n27680);
   U247 : BUF_X1 port map( A => n27682, Z => n27679);
   U248 : BUF_X1 port map( A => n27675, Z => n27673);
   U249 : BUF_X1 port map( A => n27675, Z => n27672);
   U250 : BUF_X1 port map( A => n27668, Z => n27666);
   U251 : BUF_X1 port map( A => n27668, Z => n27665);
   U252 : BUF_X1 port map( A => n27661, Z => n27659);
   U253 : BUF_X1 port map( A => n27661, Z => n27658);
   U254 : BUF_X1 port map( A => n27654, Z => n27652);
   U255 : BUF_X1 port map( A => n27654, Z => n27651);
   U256 : BUF_X1 port map( A => n27647, Z => n27645);
   U257 : BUF_X1 port map( A => n27647, Z => n27644);
   U258 : BUF_X1 port map( A => n27640, Z => n27638);
   U259 : BUF_X1 port map( A => n27640, Z => n27637);
   U260 : BUF_X1 port map( A => n27633, Z => n27631);
   U261 : BUF_X1 port map( A => n27633, Z => n27630);
   U262 : BUF_X1 port map( A => n27626, Z => n27624);
   U263 : BUF_X1 port map( A => n27626, Z => n27623);
   U264 : BUF_X1 port map( A => n27619, Z => n27617);
   U265 : BUF_X1 port map( A => n27619, Z => n27616);
   U266 : BUF_X1 port map( A => n27612, Z => n27610);
   U267 : BUF_X1 port map( A => n27612, Z => n27609);
   U268 : BUF_X1 port map( A => n27605, Z => n27603);
   U269 : BUF_X1 port map( A => n27605, Z => n27602);
   U270 : BUF_X1 port map( A => n27598, Z => n27596);
   U271 : BUF_X1 port map( A => n27598, Z => n27595);
   U272 : BUF_X1 port map( A => n27591, Z => n27589);
   U273 : BUF_X1 port map( A => n27591, Z => n27588);
   U274 : BUF_X1 port map( A => n27584, Z => n27582);
   U275 : BUF_X1 port map( A => n27584, Z => n27581);
   U276 : BUF_X1 port map( A => n27577, Z => n27575);
   U277 : BUF_X1 port map( A => n27577, Z => n27574);
   U278 : BUF_X1 port map( A => n27570, Z => n27568);
   U279 : BUF_X1 port map( A => n27570, Z => n27567);
   U280 : BUF_X1 port map( A => n27563, Z => n27561);
   U281 : BUF_X1 port map( A => n27563, Z => n27560);
   U282 : BUF_X1 port map( A => n27556, Z => n27554);
   U283 : BUF_X1 port map( A => n27556, Z => n27553);
   U284 : BUF_X1 port map( A => n27549, Z => n27547);
   U285 : BUF_X1 port map( A => n27549, Z => n27546);
   U286 : BUF_X1 port map( A => n27542, Z => n27540);
   U287 : BUF_X1 port map( A => n27542, Z => n27539);
   U288 : BUF_X1 port map( A => n27535, Z => n27533);
   U289 : BUF_X1 port map( A => n27535, Z => n27532);
   U290 : BUF_X1 port map( A => n27528, Z => n27526);
   U291 : BUF_X1 port map( A => n27528, Z => n27525);
   U292 : BUF_X1 port map( A => n27521, Z => n27519);
   U293 : BUF_X1 port map( A => n27521, Z => n27518);
   U294 : BUF_X1 port map( A => n27514, Z => n27512);
   U295 : BUF_X1 port map( A => n27514, Z => n27511);
   U296 : BUF_X1 port map( A => n27507, Z => n27505);
   U297 : BUF_X1 port map( A => n27507, Z => n27504);
   U298 : BUF_X1 port map( A => n27500, Z => n27498);
   U299 : BUF_X1 port map( A => n27500, Z => n27497);
   U300 : BUF_X1 port map( A => n27493, Z => n27491);
   U301 : BUF_X1 port map( A => n27493, Z => n27490);
   U302 : BUF_X1 port map( A => n27486, Z => n27484);
   U303 : BUF_X1 port map( A => n27486, Z => n27483);
   U304 : BUF_X1 port map( A => n27479, Z => n27477);
   U305 : BUF_X1 port map( A => n27479, Z => n27476);
   U306 : BUF_X1 port map( A => n27472, Z => n27470);
   U307 : BUF_X1 port map( A => n27472, Z => n27469);
   U308 : BUF_X1 port map( A => n27689, Z => n27688);
   U309 : BUF_X1 port map( A => n27682, Z => n27681);
   U310 : BUF_X1 port map( A => n27675, Z => n27674);
   U311 : BUF_X1 port map( A => n27668, Z => n27667);
   U312 : BUF_X1 port map( A => n27661, Z => n27660);
   U313 : BUF_X1 port map( A => n27654, Z => n27653);
   U314 : BUF_X1 port map( A => n27647, Z => n27646);
   U315 : BUF_X1 port map( A => n27640, Z => n27639);
   U316 : BUF_X1 port map( A => n27633, Z => n27632);
   U317 : BUF_X1 port map( A => n27626, Z => n27625);
   U318 : BUF_X1 port map( A => n27619, Z => n27618);
   U319 : BUF_X1 port map( A => n27612, Z => n27611);
   U320 : BUF_X1 port map( A => n27605, Z => n27604);
   U321 : BUF_X1 port map( A => n27598, Z => n27597);
   U322 : BUF_X1 port map( A => n27591, Z => n27590);
   U323 : BUF_X1 port map( A => n27584, Z => n27583);
   U324 : BUF_X1 port map( A => n27577, Z => n27576);
   U325 : BUF_X1 port map( A => n27570, Z => n27569);
   U326 : BUF_X1 port map( A => n27563, Z => n27562);
   U327 : BUF_X1 port map( A => n27556, Z => n27555);
   U328 : BUF_X1 port map( A => n27549, Z => n27548);
   U329 : BUF_X1 port map( A => n27542, Z => n27541);
   U330 : BUF_X1 port map( A => n27535, Z => n27534);
   U331 : BUF_X1 port map( A => n27528, Z => n27527);
   U332 : BUF_X1 port map( A => n27521, Z => n27520);
   U333 : BUF_X1 port map( A => n27514, Z => n27513);
   U334 : BUF_X1 port map( A => n27507, Z => n27506);
   U335 : BUF_X1 port map( A => n27500, Z => n27499);
   U336 : BUF_X1 port map( A => n27493, Z => n27492);
   U337 : BUF_X1 port map( A => n27486, Z => n27485);
   U338 : BUF_X1 port map( A => n27479, Z => n27478);
   U339 : BUF_X1 port map( A => n27472, Z => n27471);
   U340 : INV_X1 port map( A => n808_port, ZN => n27705);
   U341 : INV_X1 port map( A => n809_port, ZN => n27706);
   U342 : INV_X1 port map( A => n805_port, ZN => n27710);
   U343 : INV_X1 port map( A => n806_port, ZN => n27711);
   U344 : INV_X1 port map( A => n652_port, ZN => n27701);
   U345 : INV_X1 port map( A => n651_port, ZN => n27707);
   U346 : INV_X1 port map( A => n795_port, ZN => n27703);
   U347 : INV_X1 port map( A => n796_port, ZN => n27702);
   U348 : INV_X1 port map( A => n673_port, ZN => n27708);
   U349 : INV_X1 port map( A => n674_port, ZN => n27709);
   U350 : BUF_X1 port map( A => n674_port, Z => n26967);
   U351 : BUF_X1 port map( A => n674_port, Z => n26968);
   U352 : BUF_X1 port map( A => n673_port, Z => n26964);
   U353 : BUF_X1 port map( A => n673_port, Z => n26965);
   U354 : BUF_X1 port map( A => n674_port, Z => n26969);
   U355 : BUF_X1 port map( A => n673_port, Z => n26966);
   U356 : AND2_X1 port map( A1 => n1870, A2 => n1863, ZN => n1293);
   U357 : BUF_X1 port map( A => n26970, Z => n27057);
   U358 : BUF_X1 port map( A => n26970, Z => n27055);
   U359 : BUF_X1 port map( A => n26970, Z => n27056);
   U360 : BUF_X1 port map( A => n26970, Z => n27058);
   U361 : BUF_X1 port map( A => n26970, Z => n27059);
   U362 : BUF_X1 port map( A => n26971, Z => n27061);
   U363 : BUF_X1 port map( A => n26971, Z => n27060);
   U364 : BUF_X1 port map( A => n27264, Z => n27265);
   U365 : BUF_X1 port map( A => n27248, Z => n27249);
   U366 : BUF_X1 port map( A => n27232, Z => n27233);
   U367 : BUF_X1 port map( A => n27216, Z => n27217);
   U368 : BUF_X1 port map( A => n27200, Z => n27201);
   U369 : BUF_X1 port map( A => n27264, Z => n27266);
   U370 : BUF_X1 port map( A => n27248, Z => n27250);
   U371 : BUF_X1 port map( A => n27232, Z => n27234);
   U372 : BUF_X1 port map( A => n27216, Z => n27218);
   U373 : BUF_X1 port map( A => n27200, Z => n27202);
   U374 : BUF_X1 port map( A => n27224, Z => n27225);
   U375 : BUF_X1 port map( A => n27208, Z => n27209);
   U376 : BUF_X1 port map( A => n27224, Z => n27226);
   U377 : BUF_X1 port map( A => n27208, Z => n27210);
   U378 : BUF_X1 port map( A => n27260, Z => n27261);
   U379 : BUF_X1 port map( A => n27244, Z => n27245);
   U380 : BUF_X1 port map( A => n27228, Z => n27229);
   U381 : BUF_X1 port map( A => n27212, Z => n27213);
   U382 : BUF_X1 port map( A => n27196, Z => n27197);
   U383 : BUF_X1 port map( A => n27260, Z => n27262);
   U384 : BUF_X1 port map( A => n27244, Z => n27246);
   U385 : BUF_X1 port map( A => n27228, Z => n27230);
   U386 : BUF_X1 port map( A => n27212, Z => n27214);
   U387 : BUF_X1 port map( A => n27196, Z => n27198);
   U388 : BUF_X1 port map( A => n27268, Z => n27269);
   U389 : BUF_X1 port map( A => n27236, Z => n27237);
   U390 : BUF_X1 port map( A => n27268, Z => n27270);
   U391 : BUF_X1 port map( A => n27236, Z => n27238);
   U392 : BUF_X1 port map( A => n27182, Z => n27183);
   U393 : BUF_X1 port map( A => n27166, Z => n27167);
   U394 : BUF_X1 port map( A => n27150, Z => n27151);
   U395 : BUF_X1 port map( A => n27134, Z => n27135);
   U396 : BUF_X1 port map( A => n27118, Z => n27119);
   U397 : BUF_X1 port map( A => n27102, Z => n27103);
   U398 : BUF_X1 port map( A => n27086, Z => n27087);
   U399 : BUF_X1 port map( A => n27070, Z => n27071);
   U400 : BUF_X1 port map( A => n27182, Z => n27184);
   U401 : BUF_X1 port map( A => n27166, Z => n27168);
   U402 : BUF_X1 port map( A => n27150, Z => n27152);
   U403 : BUF_X1 port map( A => n27134, Z => n27136);
   U404 : BUF_X1 port map( A => n27118, Z => n27120);
   U405 : BUF_X1 port map( A => n27102, Z => n27104);
   U406 : BUF_X1 port map( A => n27086, Z => n27088);
   U407 : BUF_X1 port map( A => n27070, Z => n27072);
   U408 : BUF_X1 port map( A => n27178, Z => n27179);
   U409 : BUF_X1 port map( A => n27162, Z => n27163);
   U410 : BUF_X1 port map( A => n27146, Z => n27147);
   U411 : BUF_X1 port map( A => n27130, Z => n27131);
   U412 : BUF_X1 port map( A => n27114, Z => n27115);
   U413 : BUF_X1 port map( A => n27082, Z => n27083);
   U414 : BUF_X1 port map( A => n27066, Z => n27067);
   U415 : BUF_X1 port map( A => n27178, Z => n27180);
   U416 : BUF_X1 port map( A => n27162, Z => n27164);
   U417 : BUF_X1 port map( A => n27146, Z => n27148);
   U418 : BUF_X1 port map( A => n27130, Z => n27132);
   U419 : BUF_X1 port map( A => n27114, Z => n27116);
   U420 : BUF_X1 port map( A => n27082, Z => n27084);
   U421 : BUF_X1 port map( A => n27066, Z => n27068);
   U422 : BUF_X1 port map( A => n27272, Z => n27273);
   U423 : BUF_X1 port map( A => n27256, Z => n27257);
   U424 : BUF_X1 port map( A => n27240, Z => n27241);
   U425 : BUF_X1 port map( A => n27272, Z => n27274);
   U426 : BUF_X1 port map( A => n27256, Z => n27258);
   U427 : BUF_X1 port map( A => n27240, Z => n27242);
   U428 : BUF_X1 port map( A => n27186, Z => n27187);
   U429 : BUF_X1 port map( A => n27170, Z => n27171);
   U430 : BUF_X1 port map( A => n27154, Z => n27155);
   U431 : BUF_X1 port map( A => n27138, Z => n27139);
   U432 : BUF_X1 port map( A => n27122, Z => n27123);
   U433 : BUF_X1 port map( A => n27106, Z => n27107);
   U434 : BUF_X1 port map( A => n27090, Z => n27091);
   U435 : BUF_X1 port map( A => n27074, Z => n27075);
   U436 : BUF_X1 port map( A => n27186, Z => n27188);
   U437 : BUF_X1 port map( A => n27170, Z => n27172);
   U438 : BUF_X1 port map( A => n27154, Z => n27156);
   U439 : BUF_X1 port map( A => n27138, Z => n27140);
   U440 : BUF_X1 port map( A => n27122, Z => n27124);
   U441 : BUF_X1 port map( A => n27106, Z => n27108);
   U442 : BUF_X1 port map( A => n27090, Z => n27092);
   U443 : BUF_X1 port map( A => n27074, Z => n27076);
   U444 : BUF_X1 port map( A => n27252, Z => n27253);
   U445 : BUF_X1 port map( A => n27220, Z => n27221);
   U446 : BUF_X1 port map( A => n27204, Z => n27205);
   U447 : BUF_X1 port map( A => n27252, Z => n27254);
   U448 : BUF_X1 port map( A => n27220, Z => n27222);
   U449 : BUF_X1 port map( A => n27204, Z => n27206);
   U450 : BUF_X1 port map( A => n27174, Z => n27175);
   U451 : BUF_X1 port map( A => n27158, Z => n27159);
   U452 : BUF_X1 port map( A => n27142, Z => n27143);
   U453 : BUF_X1 port map( A => n27126, Z => n27127);
   U454 : BUF_X1 port map( A => n27110, Z => n27111);
   U455 : BUF_X1 port map( A => n27094, Z => n27095);
   U456 : BUF_X1 port map( A => n27078, Z => n27079);
   U457 : BUF_X1 port map( A => n27062, Z => n27063);
   U458 : BUF_X1 port map( A => n27174, Z => n27176);
   U459 : BUF_X1 port map( A => n27158, Z => n27160);
   U460 : BUF_X1 port map( A => n27142, Z => n27144);
   U461 : BUF_X1 port map( A => n27126, Z => n27128);
   U462 : BUF_X1 port map( A => n27110, Z => n27112);
   U463 : BUF_X1 port map( A => n27094, Z => n27096);
   U464 : BUF_X1 port map( A => n27078, Z => n27080);
   U465 : BUF_X1 port map( A => n27062, Z => n27064);
   U466 : BUF_X1 port map( A => n27268, Z => n27271);
   U467 : BUF_X1 port map( A => n27236, Z => n27239);
   U468 : BUF_X1 port map( A => n27182, Z => n27185);
   U469 : BUF_X1 port map( A => n27166, Z => n27169);
   U470 : BUF_X1 port map( A => n27150, Z => n27153);
   U471 : BUF_X1 port map( A => n27134, Z => n27137);
   U472 : BUF_X1 port map( A => n27118, Z => n27121);
   U473 : BUF_X1 port map( A => n27102, Z => n27105);
   U474 : BUF_X1 port map( A => n27086, Z => n27089);
   U475 : BUF_X1 port map( A => n27070, Z => n27073);
   U476 : BUF_X1 port map( A => n26962, Z => n27195);
   U477 : BUF_X1 port map( A => n26963, Z => n27192);
   U478 : BUF_X1 port map( A => n27178, Z => n27181);
   U479 : BUF_X1 port map( A => n27162, Z => n27165);
   U480 : BUF_X1 port map( A => n27146, Z => n27149);
   U481 : BUF_X1 port map( A => n27130, Z => n27133);
   U482 : BUF_X1 port map( A => n27114, Z => n27117);
   U483 : BUF_X1 port map( A => n27082, Z => n27085);
   U484 : BUF_X1 port map( A => n27066, Z => n27069);
   U485 : BUF_X1 port map( A => n27272, Z => n27275);
   U486 : BUF_X1 port map( A => n27256, Z => n27259);
   U487 : BUF_X1 port map( A => n27240, Z => n27243);
   U488 : BUF_X1 port map( A => n27186, Z => n27189);
   U489 : BUF_X1 port map( A => n27170, Z => n27173);
   U490 : BUF_X1 port map( A => n27154, Z => n27157);
   U491 : BUF_X1 port map( A => n27138, Z => n27141);
   U492 : BUF_X1 port map( A => n27122, Z => n27125);
   U493 : BUF_X1 port map( A => n27106, Z => n27109);
   U494 : BUF_X1 port map( A => n27090, Z => n27093);
   U495 : BUF_X1 port map( A => n27074, Z => n27077);
   U496 : BUF_X1 port map( A => n27252, Z => n27255);
   U497 : BUF_X1 port map( A => n27220, Z => n27223);
   U498 : BUF_X1 port map( A => n27204, Z => n27207);
   U499 : BUF_X1 port map( A => n27174, Z => n27177);
   U500 : BUF_X1 port map( A => n27158, Z => n27161);
   U501 : BUF_X1 port map( A => n27142, Z => n27145);
   U502 : BUF_X1 port map( A => n27126, Z => n27129);
   U503 : BUF_X1 port map( A => n27110, Z => n27113);
   U504 : BUF_X1 port map( A => n27094, Z => n27097);
   U505 : BUF_X1 port map( A => n27078, Z => n27081);
   U506 : BUF_X1 port map( A => n27062, Z => n27065);
   U507 : BUF_X1 port map( A => n27264, Z => n27267);
   U508 : BUF_X1 port map( A => n27248, Z => n27251);
   U509 : BUF_X1 port map( A => n27232, Z => n27235);
   U510 : BUF_X1 port map( A => n27216, Z => n27219);
   U511 : BUF_X1 port map( A => n27200, Z => n27203);
   U512 : BUF_X1 port map( A => n27224, Z => n27227);
   U513 : BUF_X1 port map( A => n27208, Z => n27211);
   U514 : BUF_X1 port map( A => n27260, Z => n27263);
   U515 : BUF_X1 port map( A => n27244, Z => n27247);
   U516 : BUF_X1 port map( A => n27228, Z => n27231);
   U517 : BUF_X1 port map( A => n27212, Z => n27215);
   U518 : BUF_X1 port map( A => n27196, Z => n27199);
   U519 : BUF_X1 port map( A => n27466, Z => n27464);
   U520 : BUF_X1 port map( A => n27460, Z => n27458);
   U521 : BUF_X1 port map( A => n27454, Z => n27452);
   U522 : BUF_X1 port map( A => n27448, Z => n27446);
   U523 : BUF_X1 port map( A => n27442, Z => n27440);
   U524 : BUF_X1 port map( A => n27280, Z => n27278);
   U525 : BUF_X1 port map( A => n27370, Z => n27368);
   U526 : BUF_X1 port map( A => n27364, Z => n27362);
   U527 : BUF_X1 port map( A => n27358, Z => n27356);
   U528 : BUF_X1 port map( A => n27352, Z => n27350);
   U529 : BUF_X1 port map( A => n27346, Z => n27344);
   U530 : BUF_X1 port map( A => n27340, Z => n27338);
   U531 : BUF_X1 port map( A => n27334, Z => n27332);
   U532 : BUF_X1 port map( A => n27328, Z => n27326);
   U533 : BUF_X1 port map( A => n27322, Z => n27320);
   U534 : BUF_X1 port map( A => n27316, Z => n27314);
   U535 : BUF_X1 port map( A => n27310, Z => n27308);
   U536 : BUF_X1 port map( A => n27304, Z => n27302);
   U537 : BUF_X1 port map( A => n27298, Z => n27296);
   U538 : BUF_X1 port map( A => n27292, Z => n27290);
   U539 : BUF_X1 port map( A => n27286, Z => n27284);
   U540 : BUF_X1 port map( A => n27436, Z => n27434);
   U541 : BUF_X1 port map( A => n27430, Z => n27428);
   U542 : BUF_X1 port map( A => n27424, Z => n27422);
   U543 : BUF_X1 port map( A => n27418, Z => n27416);
   U544 : BUF_X1 port map( A => n27412, Z => n27410);
   U545 : BUF_X1 port map( A => n27406, Z => n27404);
   U546 : BUF_X1 port map( A => n27400, Z => n27398);
   U547 : BUF_X1 port map( A => n27394, Z => n27392);
   U548 : BUF_X1 port map( A => n27388, Z => n27386);
   U549 : BUF_X1 port map( A => n27382, Z => n27380);
   U550 : BUF_X1 port map( A => n27376, Z => n27374);
   U551 : BUF_X1 port map( A => n27466, Z => n27463);
   U552 : BUF_X1 port map( A => n27460, Z => n27457);
   U553 : BUF_X1 port map( A => n27454, Z => n27451);
   U554 : BUF_X1 port map( A => n27448, Z => n27445);
   U555 : BUF_X1 port map( A => n27442, Z => n27439);
   U556 : BUF_X1 port map( A => n27280, Z => n27277);
   U557 : BUF_X1 port map( A => n27370, Z => n27367);
   U558 : BUF_X1 port map( A => n27364, Z => n27361);
   U559 : BUF_X1 port map( A => n27358, Z => n27355);
   U560 : BUF_X1 port map( A => n27352, Z => n27349);
   U561 : BUF_X1 port map( A => n27346, Z => n27343);
   U562 : BUF_X1 port map( A => n27340, Z => n27337);
   U563 : BUF_X1 port map( A => n27334, Z => n27331);
   U564 : BUF_X1 port map( A => n27328, Z => n27325);
   U565 : BUF_X1 port map( A => n27322, Z => n27319);
   U566 : BUF_X1 port map( A => n27316, Z => n27313);
   U567 : BUF_X1 port map( A => n27310, Z => n27307);
   U568 : BUF_X1 port map( A => n27304, Z => n27301);
   U569 : BUF_X1 port map( A => n27298, Z => n27295);
   U570 : BUF_X1 port map( A => n27292, Z => n27289);
   U571 : BUF_X1 port map( A => n27286, Z => n27283);
   U572 : BUF_X1 port map( A => n27436, Z => n27433);
   U573 : BUF_X1 port map( A => n27430, Z => n27427);
   U574 : BUF_X1 port map( A => n27424, Z => n27421);
   U575 : BUF_X1 port map( A => n27418, Z => n27415);
   U576 : BUF_X1 port map( A => n27412, Z => n27409);
   U577 : BUF_X1 port map( A => n27406, Z => n27403);
   U578 : BUF_X1 port map( A => n27400, Z => n27397);
   U579 : BUF_X1 port map( A => n27394, Z => n27391);
   U580 : BUF_X1 port map( A => n27388, Z => n27385);
   U581 : BUF_X1 port map( A => n27382, Z => n27379);
   U582 : BUF_X1 port map( A => n27376, Z => n27373);
   U583 : BUF_X1 port map( A => n27690, Z => n27685);
   U584 : BUF_X1 port map( A => n27691, Z => n27690);
   U585 : BUF_X1 port map( A => n27683, Z => n27678);
   U586 : BUF_X1 port map( A => n27684, Z => n27683);
   U587 : BUF_X1 port map( A => n27676, Z => n27671);
   U588 : BUF_X1 port map( A => n27677, Z => n27676);
   U589 : BUF_X1 port map( A => n27669, Z => n27664);
   U590 : BUF_X1 port map( A => n27670, Z => n27669);
   U591 : BUF_X1 port map( A => n27662, Z => n27657);
   U592 : BUF_X1 port map( A => n27663, Z => n27662);
   U593 : BUF_X1 port map( A => n27655, Z => n27650);
   U594 : BUF_X1 port map( A => n27656, Z => n27655);
   U595 : BUF_X1 port map( A => n27648, Z => n27643);
   U596 : BUF_X1 port map( A => n27649, Z => n27648);
   U597 : BUF_X1 port map( A => n27641, Z => n27636);
   U598 : BUF_X1 port map( A => n27642, Z => n27641);
   U599 : BUF_X1 port map( A => n27634, Z => n27629);
   U600 : BUF_X1 port map( A => n27635, Z => n27634);
   U601 : BUF_X1 port map( A => n27627, Z => n27622);
   U602 : BUF_X1 port map( A => n27628, Z => n27627);
   U603 : BUF_X1 port map( A => n27620, Z => n27615);
   U604 : BUF_X1 port map( A => n27621, Z => n27620);
   U605 : BUF_X1 port map( A => n27613, Z => n27608);
   U606 : BUF_X1 port map( A => n27614, Z => n27613);
   U607 : BUF_X1 port map( A => n27606, Z => n27601);
   U608 : BUF_X1 port map( A => n27607, Z => n27606);
   U609 : BUF_X1 port map( A => n27599, Z => n27594);
   U610 : BUF_X1 port map( A => n27600, Z => n27599);
   U611 : BUF_X1 port map( A => n27592, Z => n27587);
   U612 : BUF_X1 port map( A => n27593, Z => n27592);
   U613 : BUF_X1 port map( A => n27585, Z => n27580);
   U614 : BUF_X1 port map( A => n27586, Z => n27585);
   U615 : BUF_X1 port map( A => n27578, Z => n27573);
   U616 : BUF_X1 port map( A => n27579, Z => n27578);
   U617 : BUF_X1 port map( A => n27571, Z => n27566);
   U618 : BUF_X1 port map( A => n27572, Z => n27571);
   U619 : BUF_X1 port map( A => n27564, Z => n27559);
   U620 : BUF_X1 port map( A => n27565, Z => n27564);
   U621 : BUF_X1 port map( A => n27557, Z => n27552);
   U622 : BUF_X1 port map( A => n27558, Z => n27557);
   U623 : BUF_X1 port map( A => n27550, Z => n27545);
   U624 : BUF_X1 port map( A => n27551, Z => n27550);
   U625 : BUF_X1 port map( A => n27543, Z => n27538);
   U626 : BUF_X1 port map( A => n27544, Z => n27543);
   U627 : BUF_X1 port map( A => n27536, Z => n27531);
   U628 : BUF_X1 port map( A => n27537, Z => n27536);
   U629 : BUF_X1 port map( A => n27529, Z => n27524);
   U630 : BUF_X1 port map( A => n27530, Z => n27529);
   U631 : BUF_X1 port map( A => n27522, Z => n27517);
   U632 : BUF_X1 port map( A => n27523, Z => n27522);
   U633 : BUF_X1 port map( A => n27515, Z => n27510);
   U634 : BUF_X1 port map( A => n27516, Z => n27515);
   U635 : BUF_X1 port map( A => n27508, Z => n27503);
   U636 : BUF_X1 port map( A => n27509, Z => n27508);
   U637 : BUF_X1 port map( A => n27501, Z => n27496);
   U638 : BUF_X1 port map( A => n27502, Z => n27501);
   U639 : BUF_X1 port map( A => n27494, Z => n27489);
   U640 : BUF_X1 port map( A => n27495, Z => n27494);
   U641 : BUF_X1 port map( A => n27487, Z => n27482);
   U642 : BUF_X1 port map( A => n27488, Z => n27487);
   U643 : BUF_X1 port map( A => n27480, Z => n27475);
   U644 : BUF_X1 port map( A => n27481, Z => n27480);
   U645 : BUF_X1 port map( A => n27473, Z => n27468);
   U646 : BUF_X1 port map( A => n27474, Z => n27473);
   U647 : BUF_X1 port map( A => n27466, Z => n27465);
   U648 : BUF_X1 port map( A => n27460, Z => n27459);
   U649 : BUF_X1 port map( A => n27454, Z => n27453);
   U650 : BUF_X1 port map( A => n27448, Z => n27447);
   U651 : BUF_X1 port map( A => n27442, Z => n27441);
   U652 : BUF_X1 port map( A => n27280, Z => n27279);
   U653 : BUF_X1 port map( A => n27370, Z => n27369);
   U654 : BUF_X1 port map( A => n27364, Z => n27363);
   U655 : BUF_X1 port map( A => n27358, Z => n27357);
   U656 : BUF_X1 port map( A => n27352, Z => n27351);
   U657 : BUF_X1 port map( A => n27346, Z => n27345);
   U658 : BUF_X1 port map( A => n27340, Z => n27339);
   U659 : BUF_X1 port map( A => n27334, Z => n27333);
   U660 : BUF_X1 port map( A => n27328, Z => n27327);
   U661 : BUF_X1 port map( A => n27322, Z => n27321);
   U662 : BUF_X1 port map( A => n27316, Z => n27315);
   U663 : BUF_X1 port map( A => n27310, Z => n27309);
   U664 : BUF_X1 port map( A => n27304, Z => n27303);
   U665 : BUF_X1 port map( A => n27298, Z => n27297);
   U666 : BUF_X1 port map( A => n27292, Z => n27291);
   U667 : BUF_X1 port map( A => n27286, Z => n27285);
   U668 : BUF_X1 port map( A => n27436, Z => n27435);
   U669 : BUF_X1 port map( A => n27430, Z => n27429);
   U670 : BUF_X1 port map( A => n27424, Z => n27423);
   U671 : BUF_X1 port map( A => n27418, Z => n27417);
   U672 : BUF_X1 port map( A => n27412, Z => n27411);
   U673 : BUF_X1 port map( A => n27406, Z => n27405);
   U674 : BUF_X1 port map( A => n27400, Z => n27399);
   U675 : BUF_X1 port map( A => n27394, Z => n27393);
   U676 : BUF_X1 port map( A => n27388, Z => n27387);
   U677 : BUF_X1 port map( A => n27382, Z => n27381);
   U678 : BUF_X1 port map( A => n27376, Z => n27375);
   U679 : NAND2_X1 port map( A1 => n1232, A2 => n1243, ZN => n796_port);
   U680 : NAND2_X1 port map( A1 => n1236, A2 => n1240, ZN => n795_port);
   U681 : NAND2_X1 port map( A1 => n1243, A2 => n1240, ZN => n652_port);
   U682 : NAND2_X1 port map( A1 => n1235, A2 => n1240, ZN => n651_port);
   U683 : NOR2_X1 port map( A1 => n27719, A2 => n27718, ZN => n1870);
   U684 : NAND2_X1 port map( A1 => n1250, A2 => n1233, ZN => n806_port);
   U685 : NAND2_X1 port map( A1 => n1251, A2 => n1233, ZN => n805_port);
   U686 : NOR3_X1 port map( A1 => n27712, A2 => n27704, A3 => n27713, ZN => 
                           n1241);
   U687 : NAND2_X1 port map( A1 => n1250, A2 => n1235, ZN => n809_port);
   U688 : NAND2_X1 port map( A1 => n1251, A2 => n1235, ZN => n808_port);
   U689 : NOR3_X1 port map( A1 => n27716, A2 => n27715, A3 => n27717, ZN => 
                           n1863);
   U690 : NAND2_X1 port map( A1 => n1251, A2 => n1234, ZN => n674_port);
   U691 : NAND2_X1 port map( A1 => n1250, A2 => n1234, ZN => n673_port);
   U692 : AND2_X1 port map( A1 => n1250, A2 => n1236, ZN => n26962);
   U693 : AND2_X1 port map( A1 => n1251, A2 => n1236, ZN => n26963);
   U694 : NAND2_X1 port map( A1 => n955_port, A2 => n956_port, ZN => out2(23));
   U695 : NOR4_X1 port map( A1 => n965_port, A2 => n966_port, A3 => n967_port, 
                           A4 => n968_port, ZN => n955_port);
   U696 : NOR4_X1 port map( A1 => n957_port, A2 => n958_port, A3 => n959_port, 
                           A4 => n960_port, ZN => n956_port);
   U697 : OAI221_X1 port map( B1 => n27210, B2 => n26655, C1 => n27206, C2 => 
                           n26382, A => n970_port, ZN => n967_port);
   U698 : NAND2_X1 port map( A1 => n937_port, A2 => n938_port, ZN => out2(24));
   U699 : NOR4_X1 port map( A1 => n947_port, A2 => n948_port, A3 => n949_port, 
                           A4 => n950_port, ZN => n937_port);
   U700 : NOR4_X1 port map( A1 => n939_port, A2 => n940_port, A3 => n941_port, 
                           A4 => n942_port, ZN => n938_port);
   U701 : OAI221_X1 port map( B1 => n27210, B2 => n26656, C1 => n27206, C2 => 
                           n26383, A => n952_port, ZN => n949_port);
   U702 : NAND2_X1 port map( A1 => n919_port, A2 => n920_port, ZN => out2(25));
   U703 : NOR4_X1 port map( A1 => n929_port, A2 => n930_port, A3 => n931_port, 
                           A4 => n932_port, ZN => n919_port);
   U704 : NOR4_X1 port map( A1 => n921_port, A2 => n922_port, A3 => n923_port, 
                           A4 => n924_port, ZN => n920_port);
   U705 : OAI221_X1 port map( B1 => n27210, B2 => n26657, C1 => n27206, C2 => 
                           n26384, A => n934_port, ZN => n931_port);
   U706 : NAND2_X1 port map( A1 => n901_port, A2 => n902_port, ZN => out2(26));
   U707 : NOR4_X1 port map( A1 => n911_port, A2 => n912_port, A3 => n913_port, 
                           A4 => n914_port, ZN => n901_port);
   U708 : NOR4_X1 port map( A1 => n903_port, A2 => n904_port, A3 => n905_port, 
                           A4 => n906_port, ZN => n902_port);
   U709 : OAI221_X1 port map( B1 => n27210, B2 => n26658, C1 => n27206, C2 => 
                           n26385, A => n916_port, ZN => n913_port);
   U710 : NAND2_X1 port map( A1 => n883_port, A2 => n884_port, ZN => out2(27));
   U711 : NOR4_X1 port map( A1 => n893_port, A2 => n894_port, A3 => n895_port, 
                           A4 => n896_port, ZN => n883_port);
   U712 : NOR4_X1 port map( A1 => n885_port, A2 => n886_port, A3 => n887_port, 
                           A4 => n888_port, ZN => n884_port);
   U713 : OAI221_X1 port map( B1 => n27210, B2 => n26659, C1 => n27206, C2 => 
                           n26386, A => n898_port, ZN => n895_port);
   U714 : NAND2_X1 port map( A1 => n865_port, A2 => n866_port, ZN => out2(28));
   U715 : NOR4_X1 port map( A1 => n875_port, A2 => n876_port, A3 => n877_port, 
                           A4 => n878_port, ZN => n865_port);
   U716 : NOR4_X1 port map( A1 => n867_port, A2 => n868_port, A3 => n869_port, 
                           A4 => n870_port, ZN => n866_port);
   U717 : OAI221_X1 port map( B1 => n27210, B2 => n26660, C1 => n27206, C2 => 
                           n26387, A => n880_port, ZN => n877_port);
   U718 : NAND2_X1 port map( A1 => n847_port, A2 => n848_port, ZN => out2(29));
   U719 : NOR4_X1 port map( A1 => n857_port, A2 => n858_port, A3 => n859_port, 
                           A4 => n860_port, ZN => n847_port);
   U720 : NOR4_X1 port map( A1 => n849_port, A2 => n850_port, A3 => n851_port, 
                           A4 => n852_port, ZN => n848_port);
   U721 : OAI221_X1 port map( B1 => n27210, B2 => n26661, C1 => n27206, C2 => 
                           n26388, A => n862_port, ZN => n859_port);
   U722 : NAND2_X1 port map( A1 => n811_port, A2 => n812_port, ZN => out2(30));
   U723 : NOR4_X1 port map( A1 => n821_port, A2 => n822_port, A3 => n823_port, 
                           A4 => n824_port, ZN => n811_port);
   U724 : NOR4_X1 port map( A1 => n813_port, A2 => n814_port, A3 => n815_port, 
                           A4 => n816_port, ZN => n812_port);
   U725 : OAI221_X1 port map( B1 => n27210, B2 => n26662, C1 => n27207, C2 => 
                           n26389, A => n826_port, ZN => n823_port);
   U726 : NAND2_X1 port map( A1 => n787_port, A2 => n788_port, ZN => out2(31));
   U727 : NOR4_X1 port map( A1 => n799_port, A2 => n800_port, A3 => n801_port, 
                           A4 => n802_port, ZN => n787_port);
   U728 : NOR4_X1 port map( A1 => n789_port, A2 => n790_port, A3 => n791_port, 
                           A4 => n792_port, ZN => n788_port);
   U729 : OAI221_X1 port map( B1 => n27211, B2 => n26663, C1 => n27207, C2 => 
                           n26390, A => n804_port, ZN => n801_port);
   U730 : NAND2_X1 port map( A1 => n1845, A2 => n1846, ZN => out1(0));
   U731 : NOR4_X1 port map( A1 => n1865, A2 => n1866, A3 => n1867, A4 => n1868,
                           ZN => n1845);
   U732 : NOR4_X1 port map( A1 => n1847, A2 => n1848, A3 => n1849, A4 => n1850,
                           ZN => n1846);
   U733 : OAI221_X1 port map( B1 => n26498, B2 => n27075, C1 => n26814, C2 => 
                           n27071, A => n1874, ZN => n1865);
   U734 : NAND2_X1 port map( A1 => n1647, A2 => n1648, ZN => out1(1));
   U735 : NOR4_X1 port map( A1 => n1657, A2 => n1658, A3 => n1659, A4 => n1660,
                           ZN => n1647);
   U736 : NOR4_X1 port map( A1 => n1649, A2 => n1650, A3 => n1651, A4 => n1652,
                           ZN => n1648);
   U737 : OAI221_X1 port map( B1 => n26499, B2 => n27076, C1 => n26815, C2 => 
                           n27072, A => n1664, ZN => n1657);
   U738 : NAND2_X1 port map( A1 => n1449, A2 => n1450, ZN => out1(2));
   U739 : NOR4_X1 port map( A1 => n1459, A2 => n1460, A3 => n1461, A4 => n1462,
                           ZN => n1449);
   U740 : NOR4_X1 port map( A1 => n1451, A2 => n1452, A3 => n1453, A4 => n1454,
                           ZN => n1450);
   U741 : OAI221_X1 port map( B1 => n26500, B2 => n27077, C1 => n26816, C2 => 
                           n27073, A => n1466, ZN => n1459);
   U742 : NAND2_X1 port map( A1 => n1395, A2 => n1396, ZN => out1(3));
   U743 : NOR4_X1 port map( A1 => n1405, A2 => n1406, A3 => n1407, A4 => n1408,
                           ZN => n1395);
   U744 : NOR4_X1 port map( A1 => n1397, A2 => n1398, A3 => n1399, A4 => n1400,
                           ZN => n1396);
   U745 : OAI221_X1 port map( B1 => n26501, B2 => n27077, C1 => n26817, C2 => 
                           n27073, A => n1412, ZN => n1405);
   U746 : NAND2_X1 port map( A1 => n1377, A2 => n1378, ZN => out1(4));
   U747 : NOR4_X1 port map( A1 => n1387, A2 => n1388, A3 => n1389, A4 => n1390,
                           ZN => n1377);
   U748 : NOR4_X1 port map( A1 => n1379, A2 => n1380, A3 => n1381, A4 => n1382,
                           ZN => n1378);
   U749 : OAI221_X1 port map( B1 => n26502, B2 => n27077, C1 => n26818, C2 => 
                           n27073, A => n1394, ZN => n1387);
   U750 : NAND2_X1 port map( A1 => n1359, A2 => n1360, ZN => out1(5));
   U751 : NOR4_X1 port map( A1 => n1369, A2 => n1370, A3 => n1371, A4 => n1372,
                           ZN => n1359);
   U752 : NOR4_X1 port map( A1 => n1361, A2 => n1362, A3 => n1363, A4 => n1364,
                           ZN => n1360);
   U753 : OAI221_X1 port map( B1 => n26503, B2 => n27077, C1 => n26819, C2 => 
                           n27073, A => n1376, ZN => n1369);
   U754 : NAND2_X1 port map( A1 => n1341, A2 => n1342, ZN => out1(6));
   U755 : NOR4_X1 port map( A1 => n1351, A2 => n1352, A3 => n1353, A4 => n1354,
                           ZN => n1341);
   U756 : NOR4_X1 port map( A1 => n1343, A2 => n1344, A3 => n1345, A4 => n1346,
                           ZN => n1342);
   U757 : OAI221_X1 port map( B1 => n26504, B2 => n27077, C1 => n26820, C2 => 
                           n27073, A => n1358, ZN => n1351);
   U758 : NAND2_X1 port map( A1 => n1323, A2 => n1324, ZN => out1(7));
   U759 : NOR4_X1 port map( A1 => n1333, A2 => n1334, A3 => n1335, A4 => n1336,
                           ZN => n1323);
   U760 : NOR4_X1 port map( A1 => n1325, A2 => n1326, A3 => n1327, A4 => n1328,
                           ZN => n1324);
   U761 : OAI221_X1 port map( B1 => n26505, B2 => n27077, C1 => n26821, C2 => 
                           n27073, A => n1340, ZN => n1333);
   U762 : NAND2_X1 port map( A1 => n1305, A2 => n1306, ZN => out1(8));
   U763 : NOR4_X1 port map( A1 => n1315, A2 => n1316, A3 => n1317, A4 => n1318,
                           ZN => n1305);
   U764 : NOR4_X1 port map( A1 => n1307, A2 => n1308, A3 => n1309, A4 => n1310,
                           ZN => n1306);
   U765 : OAI221_X1 port map( B1 => n26506, B2 => n27077, C1 => n26822, C2 => 
                           n27073, A => n1322, ZN => n1315);
   U766 : NAND2_X1 port map( A1 => n1255, A2 => n1256, ZN => out1(9));
   U767 : NOR4_X1 port map( A1 => n1281, A2 => n1282, A3 => n1283, A4 => n1284,
                           ZN => n1255);
   U768 : NOR4_X1 port map( A1 => n1257, A2 => n1258, A3 => n1259, A4 => n1260,
                           ZN => n1256);
   U769 : OAI221_X1 port map( B1 => n26507, B2 => n27077, C1 => n26823, C2 => 
                           n27073, A => n1302, ZN => n1281);
   U770 : NAND2_X1 port map( A1 => n1827, A2 => n1828, ZN => out1(10));
   U771 : NOR4_X1 port map( A1 => n1837, A2 => n1838, A3 => n1839, A4 => n1840,
                           ZN => n1827);
   U772 : NOR4_X1 port map( A1 => n1829, A2 => n1830, A3 => n1831, A4 => n1832,
                           ZN => n1828);
   U773 : OAI221_X1 port map( B1 => n26508, B2 => n27075, C1 => n26824, C2 => 
                           n27071, A => n1844, ZN => n1837);
   U774 : NAND2_X1 port map( A1 => n1809, A2 => n1810, ZN => out1(11));
   U775 : NOR4_X1 port map( A1 => n1819, A2 => n1820, A3 => n1821, A4 => n1822,
                           ZN => n1809);
   U776 : NOR4_X1 port map( A1 => n1811, A2 => n1812, A3 => n1813, A4 => n1814,
                           ZN => n1810);
   U777 : OAI221_X1 port map( B1 => n26509, B2 => n27075, C1 => n26825, C2 => 
                           n27071, A => n1826, ZN => n1819);
   U778 : NAND2_X1 port map( A1 => n1791, A2 => n1792, ZN => out1(12));
   U779 : NOR4_X1 port map( A1 => n1801, A2 => n1802, A3 => n1803, A4 => n1804,
                           ZN => n1791);
   U780 : NOR4_X1 port map( A1 => n1793, A2 => n1794, A3 => n1795, A4 => n1796,
                           ZN => n1792);
   U781 : OAI221_X1 port map( B1 => n26510, B2 => n27075, C1 => n26826, C2 => 
                           n27071, A => n1808, ZN => n1801);
   U782 : NAND2_X1 port map( A1 => n1773, A2 => n1774, ZN => out1(13));
   U783 : NOR4_X1 port map( A1 => n1783, A2 => n1784, A3 => n1785, A4 => n1786,
                           ZN => n1773);
   U784 : NOR4_X1 port map( A1 => n1775, A2 => n1776, A3 => n1777, A4 => n1778,
                           ZN => n1774);
   U785 : OAI221_X1 port map( B1 => n26511, B2 => n27075, C1 => n26827, C2 => 
                           n27071, A => n1790, ZN => n1783);
   U786 : NAND2_X1 port map( A1 => n1755, A2 => n1756, ZN => out1(14));
   U787 : NOR4_X1 port map( A1 => n1765, A2 => n1766, A3 => n1767, A4 => n1768,
                           ZN => n1755);
   U788 : NOR4_X1 port map( A1 => n1757, A2 => n1758, A3 => n1759, A4 => n1760,
                           ZN => n1756);
   U789 : OAI221_X1 port map( B1 => n26512, B2 => n27075, C1 => n26828, C2 => 
                           n27071, A => n1772, ZN => n1765);
   U790 : NAND2_X1 port map( A1 => n1737, A2 => n1738, ZN => out1(15));
   U791 : NOR4_X1 port map( A1 => n1747, A2 => n1748, A3 => n1749, A4 => n1750,
                           ZN => n1737);
   U792 : NOR4_X1 port map( A1 => n1739, A2 => n1740, A3 => n1741, A4 => n1742,
                           ZN => n1738);
   U793 : OAI221_X1 port map( B1 => n26513, B2 => n27075, C1 => n26829, C2 => 
                           n27071, A => n1754, ZN => n1747);
   U794 : NAND2_X1 port map( A1 => n1719, A2 => n1720, ZN => out1(16));
   U795 : NOR4_X1 port map( A1 => n1729, A2 => n1730, A3 => n1731, A4 => n1732,
                           ZN => n1719);
   U796 : NOR4_X1 port map( A1 => n1721, A2 => n1722, A3 => n1723, A4 => n1724,
                           ZN => n1720);
   U797 : OAI221_X1 port map( B1 => n26514, B2 => n27075, C1 => n26830, C2 => 
                           n27071, A => n1736, ZN => n1729);
   U798 : NAND2_X1 port map( A1 => n1701, A2 => n1702, ZN => out1(17));
   U799 : NOR4_X1 port map( A1 => n1711, A2 => n1712, A3 => n1713, A4 => n1714,
                           ZN => n1701);
   U800 : NOR4_X1 port map( A1 => n1703, A2 => n1704, A3 => n1705, A4 => n1706,
                           ZN => n1702);
   U801 : OAI221_X1 port map( B1 => n26515, B2 => n27075, C1 => n26831, C2 => 
                           n27071, A => n1718, ZN => n1711);
   U802 : NAND2_X1 port map( A1 => n1683, A2 => n1684, ZN => out1(18));
   U803 : NOR4_X1 port map( A1 => n1693, A2 => n1694, A3 => n1695, A4 => n1696,
                           ZN => n1683);
   U804 : NOR4_X1 port map( A1 => n1685, A2 => n1686, A3 => n1687, A4 => n1688,
                           ZN => n1684);
   U805 : OAI221_X1 port map( B1 => n26516, B2 => n27075, C1 => n26832, C2 => 
                           n27071, A => n1700, ZN => n1693);
   U806 : NAND2_X1 port map( A1 => n1665, A2 => n1666, ZN => out1(19));
   U807 : NOR4_X1 port map( A1 => n1675, A2 => n1676, A3 => n1677, A4 => n1678,
                           ZN => n1665);
   U808 : NOR4_X1 port map( A1 => n1667, A2 => n1668, A3 => n1669, A4 => n1670,
                           ZN => n1666);
   U809 : OAI221_X1 port map( B1 => n26517, B2 => n27075, C1 => n26833, C2 => 
                           n27071, A => n1682, ZN => n1675);
   U810 : NAND2_X1 port map( A1 => n1629, A2 => n1630, ZN => out1(20));
   U811 : NOR4_X1 port map( A1 => n1639, A2 => n1640, A3 => n1641, A4 => n1642,
                           ZN => n1629);
   U812 : NOR4_X1 port map( A1 => n1631, A2 => n1632, A3 => n1633, A4 => n1634,
                           ZN => n1630);
   U813 : OAI221_X1 port map( B1 => n26518, B2 => n27076, C1 => n26834, C2 => 
                           n27072, A => n1646, ZN => n1639);
   U814 : NAND2_X1 port map( A1 => n1611, A2 => n1612, ZN => out1(21));
   U815 : NOR4_X1 port map( A1 => n1621, A2 => n1622, A3 => n1623, A4 => n1624,
                           ZN => n1611);
   U816 : NOR4_X1 port map( A1 => n1613, A2 => n1614, A3 => n1615, A4 => n1616,
                           ZN => n1612);
   U817 : OAI221_X1 port map( B1 => n26519, B2 => n27076, C1 => n26835, C2 => 
                           n27072, A => n1628, ZN => n1621);
   U818 : NAND2_X1 port map( A1 => n1593, A2 => n1594, ZN => out1(22));
   U819 : NOR4_X1 port map( A1 => n1603, A2 => n1604, A3 => n1605, A4 => n1606,
                           ZN => n1593);
   U820 : NOR4_X1 port map( A1 => n1595, A2 => n1596, A3 => n1597, A4 => n1598,
                           ZN => n1594);
   U821 : OAI221_X1 port map( B1 => n26520, B2 => n27076, C1 => n26836, C2 => 
                           n27072, A => n1610, ZN => n1603);
   U822 : NAND2_X1 port map( A1 => n1575, A2 => n1576, ZN => out1(23));
   U823 : NOR4_X1 port map( A1 => n1585, A2 => n1586, A3 => n1587, A4 => n1588,
                           ZN => n1575);
   U824 : NOR4_X1 port map( A1 => n1577, A2 => n1578, A3 => n1579, A4 => n1580,
                           ZN => n1576);
   U825 : OAI221_X1 port map( B1 => n26521, B2 => n27076, C1 => n26837, C2 => 
                           n27072, A => n1592, ZN => n1585);
   U826 : NAND2_X1 port map( A1 => n1557, A2 => n1558, ZN => out1(24));
   U827 : NOR4_X1 port map( A1 => n1567, A2 => n1568, A3 => n1569, A4 => n1570,
                           ZN => n1557);
   U828 : NOR4_X1 port map( A1 => n1559, A2 => n1560, A3 => n1561, A4 => n1562,
                           ZN => n1558);
   U829 : OAI221_X1 port map( B1 => n26522, B2 => n27076, C1 => n26838, C2 => 
                           n27072, A => n1574, ZN => n1567);
   U830 : NAND2_X1 port map( A1 => n1539, A2 => n1540, ZN => out1(25));
   U831 : NOR4_X1 port map( A1 => n1549, A2 => n1550, A3 => n1551, A4 => n1552,
                           ZN => n1539);
   U832 : NOR4_X1 port map( A1 => n1541, A2 => n1542, A3 => n1543, A4 => n1544,
                           ZN => n1540);
   U833 : OAI221_X1 port map( B1 => n26523, B2 => n27076, C1 => n26839, C2 => 
                           n27072, A => n1556, ZN => n1549);
   U834 : NAND2_X1 port map( A1 => n1521, A2 => n1522, ZN => out1(26));
   U835 : NOR4_X1 port map( A1 => n1531, A2 => n1532, A3 => n1533, A4 => n1534,
                           ZN => n1521);
   U836 : NOR4_X1 port map( A1 => n1523, A2 => n1524, A3 => n1525, A4 => n1526,
                           ZN => n1522);
   U837 : OAI221_X1 port map( B1 => n26524, B2 => n27076, C1 => n26840, C2 => 
                           n27072, A => n1538, ZN => n1531);
   U838 : NAND2_X1 port map( A1 => n1503, A2 => n1504, ZN => out1(27));
   U839 : NOR4_X1 port map( A1 => n1513, A2 => n1514, A3 => n1515, A4 => n1516,
                           ZN => n1503);
   U840 : NOR4_X1 port map( A1 => n1505, A2 => n1506, A3 => n1507, A4 => n1508,
                           ZN => n1504);
   U841 : OAI221_X1 port map( B1 => n26525, B2 => n27076, C1 => n26841, C2 => 
                           n27072, A => n1520, ZN => n1513);
   U842 : NAND2_X1 port map( A1 => n1485, A2 => n1486, ZN => out1(28));
   U843 : NOR4_X1 port map( A1 => n1495, A2 => n1496, A3 => n1497, A4 => n1498,
                           ZN => n1485);
   U844 : NOR4_X1 port map( A1 => n1487, A2 => n1488, A3 => n1489, A4 => n1490,
                           ZN => n1486);
   U845 : OAI221_X1 port map( B1 => n26526, B2 => n27076, C1 => n26842, C2 => 
                           n27072, A => n1502, ZN => n1495);
   U846 : NAND2_X1 port map( A1 => n1467, A2 => n1468, ZN => out1(29));
   U847 : NOR4_X1 port map( A1 => n1477, A2 => n1478, A3 => n1479, A4 => n1480,
                           ZN => n1467);
   U848 : NOR4_X1 port map( A1 => n1469, A2 => n1470, A3 => n1471, A4 => n1472,
                           ZN => n1468);
   U849 : OAI221_X1 port map( B1 => n26527, B2 => n27076, C1 => n26843, C2 => 
                           n27072, A => n1484, ZN => n1477);
   U850 : NAND2_X1 port map( A1 => n1431, A2 => n1432, ZN => out1(30));
   U851 : NOR4_X1 port map( A1 => n1441, A2 => n1442, A3 => n1443, A4 => n1444,
                           ZN => n1431);
   U852 : NOR4_X1 port map( A1 => n1433, A2 => n1434, A3 => n1435, A4 => n1436,
                           ZN => n1432);
   U853 : OAI221_X1 port map( B1 => n26528, B2 => n27077, C1 => n26844, C2 => 
                           n27073, A => n1448, ZN => n1441);
   U854 : NAND2_X1 port map( A1 => n1413, A2 => n1414, ZN => out1(31));
   U855 : NOR4_X1 port map( A1 => n1423, A2 => n1424, A3 => n1425, A4 => n1426,
                           ZN => n1413);
   U856 : NOR4_X1 port map( A1 => n1415, A2 => n1416, A3 => n1417, A4 => n1418,
                           ZN => n1414);
   U857 : OAI221_X1 port map( B1 => n26529, B2 => n27077, C1 => n26845, C2 => 
                           n27073, A => n1430, ZN => n1423);
   U858 : NAND2_X1 port map( A1 => n1232, A2 => n1235, ZN => n642_port);
   U859 : NAND2_X1 port map( A1 => n1232, A2 => n1236, ZN => n641_port);
   U860 : NAND2_X1 port map( A1 => n1232, A2 => n1241, ZN => n646_port);
   U861 : NAND2_X1 port map( A1 => n1234, A2 => n1240, ZN => n647_port);
   U862 : NAND2_X1 port map( A1 => n1239, A2 => n1240, ZN => n655_port);
   U863 : NAND2_X1 port map( A1 => n1241, A2 => n1240, ZN => n654_port);
   U864 : NAND2_X1 port map( A1 => n1250, A2 => n1238, ZN => n664_port);
   U865 : NAND2_X1 port map( A1 => n1251, A2 => n1238, ZN => n663_port);
   U866 : NAND2_X1 port map( A1 => n1250, A2 => n1243, ZN => n669_port);
   U867 : NAND2_X1 port map( A1 => n1251, A2 => n1243, ZN => n668_port);
   U868 : NAND2_X1 port map( A1 => n1855, A2 => n1853, ZN => n1262);
   U869 : NAND2_X1 port map( A1 => n1855, A2 => n1854, ZN => n1261);
   U870 : NAND2_X1 port map( A1 => n1858, A2 => n1853, ZN => n1267);
   U871 : NAND2_X1 port map( A1 => n1858, A2 => n1854, ZN => n1266);
   U872 : NAND2_X1 port map( A1 => n1861, A2 => n1853, ZN => n1272);
   U873 : NAND2_X1 port map( A1 => n1861, A2 => n1854, ZN => n1271);
   U874 : NAND2_X1 port map( A1 => n1864, A2 => n1853, ZN => n1277);
   U875 : NAND2_X1 port map( A1 => n1864, A2 => n1854, ZN => n1276);
   U876 : NAND2_X1 port map( A1 => n1870, A2 => n1855, ZN => n1286);
   U877 : NAND2_X1 port map( A1 => n1870, A2 => n1852, ZN => n1285);
   U878 : NAND2_X1 port map( A1 => n1870, A2 => n1861, ZN => n1291);
   U879 : NAND2_X1 port map( A1 => n1870, A2 => n1860, ZN => n1290);
   U880 : NAND2_X1 port map( A1 => n1872, A2 => n1864, ZN => n1296);
   U881 : NAND2_X1 port map( A1 => n1872, A2 => n1855, ZN => n1295);
   U882 : NAND2_X1 port map( A1 => n1872, A2 => n1861, ZN => n1301);
   U883 : NAND2_X1 port map( A1 => n1872, A2 => n1857, ZN => n1300);
   U884 : AND2_X1 port map( A1 => n1234, A2 => n1232, ZN => n644_port);
   U885 : AND2_X1 port map( A1 => n1233, A2 => n1240, ZN => n657_port);
   U886 : AND2_X1 port map( A1 => n1238, A2 => n1240, ZN => n658_port);
   U887 : AND2_X1 port map( A1 => n1251, A2 => n1239, ZN => n666_port);
   U888 : AND2_X1 port map( A1 => n1250, A2 => n1239, ZN => n667_port);
   U889 : AND2_X1 port map( A1 => n1251, A2 => n1241, ZN => n671_port);
   U890 : AND2_X1 port map( A1 => n1250, A2 => n1241, ZN => n672_port);
   U891 : AND2_X1 port map( A1 => n1853, A2 => n1863, ZN => n1280);
   U892 : AND2_X1 port map( A1 => n1870, A2 => n1858, ZN => n1288);
   U893 : AND2_X1 port map( A1 => n1870, A2 => n1857, ZN => n1289);
   U894 : AND2_X1 port map( A1 => n1872, A2 => n1858, ZN => n1294);
   U895 : AND2_X1 port map( A1 => n1872, A2 => n1852, ZN => n1298);
   U896 : AND2_X1 port map( A1 => n1870, A2 => n1864, ZN => n1299);
   U897 : AND2_X1 port map( A1 => n1872, A2 => n1863, ZN => n1303);
   U898 : AND2_X1 port map( A1 => n1872, A2 => n1860, ZN => n1304);
   U899 : AND2_X1 port map( A1 => n1232, A2 => n1233, ZN => n645_port);
   U900 : AND2_X1 port map( A1 => n1232, A2 => n1239, ZN => n649_port);
   U901 : AND2_X1 port map( A1 => n1232, A2 => n1238, ZN => n650_port);
   U902 : AND2_X1 port map( A1 => n1852, A2 => n1854, ZN => n1264);
   U903 : AND2_X1 port map( A1 => n1852, A2 => n1853, ZN => n1265);
   U904 : AND2_X1 port map( A1 => n1857, A2 => n1854, ZN => n1269);
   U905 : AND2_X1 port map( A1 => n1857, A2 => n1853, ZN => n1270);
   U906 : AND2_X1 port map( A1 => n1860, A2 => n1854, ZN => n1274);
   U907 : AND2_X1 port map( A1 => n1860, A2 => n1853, ZN => n1275);
   U908 : AND2_X1 port map( A1 => n1863, A2 => n1854, ZN => n1279);
   U909 : BUF_X1 port map( A => N2166, Z => n27691);
   U910 : OAI21_X1 port map( B1 => n1883, B2 => n1886, A => n26973, ZN => N2166
                           );
   U911 : BUF_X1 port map( A => N2199, Z => n27684);
   U912 : OAI21_X1 port map( B1 => n1882, B2 => n1886, A => n26972, ZN => N2199
                           );
   U913 : BUF_X1 port map( A => N2231, Z => n27677);
   U914 : OAI21_X1 port map( B1 => n1881, B2 => n1886, A => n26973, ZN => N2231
                           );
   U915 : BUF_X1 port map( A => N2263, Z => n27670);
   U916 : OAI21_X1 port map( B1 => n1880, B2 => n1886, A => n26973, ZN => N2263
                           );
   U917 : BUF_X1 port map( A => N2295, Z => n27663);
   U918 : OAI21_X1 port map( B1 => n1879, B2 => n1886, A => n26973, ZN => N2295
                           );
   U919 : BUF_X1 port map( A => N2327, Z => n27656);
   U920 : OAI21_X1 port map( B1 => n1878, B2 => n1886, A => n26974, ZN => N2327
                           );
   U921 : BUF_X1 port map( A => N2359, Z => n27649);
   U922 : OAI21_X1 port map( B1 => n1877, B2 => n1886, A => n26974, ZN => N2359
                           );
   U923 : BUF_X1 port map( A => N2391, Z => n27642);
   U924 : OAI21_X1 port map( B1 => n1876, B2 => n1886, A => n26974, ZN => N2391
                           );
   U925 : BUF_X1 port map( A => N2423, Z => n27635);
   U926 : OAI21_X1 port map( B1 => n1883, B2 => n1885, A => n26974, ZN => N2423
                           );
   U927 : BUF_X1 port map( A => N2455, Z => n27628);
   U928 : OAI21_X1 port map( B1 => n1882, B2 => n1885, A => n26974, ZN => N2455
                           );
   U929 : BUF_X1 port map( A => N2487, Z => n27621);
   U930 : OAI21_X1 port map( B1 => n1881, B2 => n1885, A => n26973, ZN => N2487
                           );
   U931 : BUF_X1 port map( A => N2519, Z => n27614);
   U932 : OAI21_X1 port map( B1 => n1880, B2 => n1885, A => n26974, ZN => N2519
                           );
   U933 : BUF_X1 port map( A => N2551, Z => n27607);
   U934 : OAI21_X1 port map( B1 => n1879, B2 => n1885, A => n26973, ZN => N2551
                           );
   U935 : BUF_X1 port map( A => N2583, Z => n27600);
   U936 : OAI21_X1 port map( B1 => n1878, B2 => n1885, A => n26974, ZN => N2583
                           );
   U937 : BUF_X1 port map( A => N2615, Z => n27593);
   U938 : OAI21_X1 port map( B1 => n1877, B2 => n1885, A => n26973, ZN => N2615
                           );
   U939 : BUF_X1 port map( A => N2647, Z => n27586);
   U940 : OAI21_X1 port map( B1 => n1876, B2 => n1885, A => n26974, ZN => N2647
                           );
   U941 : BUF_X1 port map( A => N2679, Z => n27579);
   U942 : OAI21_X1 port map( B1 => n1883, B2 => n1884, A => n26974, ZN => N2679
                           );
   U943 : BUF_X1 port map( A => N2711, Z => n27572);
   U944 : OAI21_X1 port map( B1 => n1882, B2 => n1884, A => n26974, ZN => N2711
                           );
   U945 : BUF_X1 port map( A => N2743, Z => n27565);
   U946 : OAI21_X1 port map( B1 => n1881, B2 => n1884, A => n26973, ZN => N2743
                           );
   U947 : BUF_X1 port map( A => N2775, Z => n27558);
   U948 : OAI21_X1 port map( B1 => n1880, B2 => n1884, A => n26973, ZN => N2775
                           );
   U949 : BUF_X1 port map( A => N2807, Z => n27551);
   U950 : OAI21_X1 port map( B1 => n1879, B2 => n1884, A => n26972, ZN => N2807
                           );
   U951 : BUF_X1 port map( A => N2839, Z => n27544);
   U952 : OAI21_X1 port map( B1 => n1878, B2 => n1884, A => n26973, ZN => N2839
                           );
   U953 : BUF_X1 port map( A => N2871, Z => n27537);
   U954 : OAI21_X1 port map( B1 => n1877, B2 => n1884, A => n26972, ZN => N2871
                           );
   U955 : BUF_X1 port map( A => N2903, Z => n27530);
   U956 : OAI21_X1 port map( B1 => n1876, B2 => n1884, A => n26972, ZN => N2903
                           );
   U957 : BUF_X1 port map( A => N2935, Z => n27523);
   U958 : OAI21_X1 port map( B1 => n1875, B2 => n1883, A => n26972, ZN => N2935
                           );
   U959 : BUF_X1 port map( A => N2967, Z => n27516);
   U960 : OAI21_X1 port map( B1 => n1875, B2 => n1882, A => n26972, ZN => N2967
                           );
   U961 : BUF_X1 port map( A => N2999, Z => n27509);
   U962 : OAI21_X1 port map( B1 => n1875, B2 => n1881, A => n26973, ZN => N2999
                           );
   U963 : BUF_X1 port map( A => N3031, Z => n27502);
   U964 : OAI21_X1 port map( B1 => n1875, B2 => n1880, A => n26972, ZN => N3031
                           );
   U965 : BUF_X1 port map( A => N3063, Z => n27495);
   U966 : OAI21_X1 port map( B1 => n1875, B2 => n1879, A => n26972, ZN => N3063
                           );
   U967 : BUF_X1 port map( A => N3095, Z => n27488);
   U968 : OAI21_X1 port map( B1 => n1875, B2 => n1878, A => n26972, ZN => N3095
                           );
   U969 : BUF_X1 port map( A => N3127, Z => n27481);
   U970 : OAI21_X1 port map( B1 => n1875, B2 => n1877, A => n26972, ZN => N3127
                           );
   U971 : BUF_X1 port map( A => N3159, Z => n27474);
   U972 : OAI21_X1 port map( B1 => n1875, B2 => n1876, A => n26972, ZN => N3159
                           );
   U973 : BUF_X1 port map( A => n27720, Z => n26971);
   U974 : BUF_X1 port map( A => n27467, Z => n27462);
   U975 : BUF_X1 port map( A => n26680, Z => n27467);
   U976 : BUF_X1 port map( A => n27461, Z => n27456);
   U977 : BUF_X1 port map( A => n26681, Z => n27461);
   U978 : BUF_X1 port map( A => n27455, Z => n27450);
   U979 : BUF_X1 port map( A => n26682, Z => n27455);
   U980 : BUF_X1 port map( A => n27449, Z => n27444);
   U981 : BUF_X1 port map( A => n26683, Z => n27449);
   U982 : BUF_X1 port map( A => n27443, Z => n27438);
   U983 : BUF_X1 port map( A => n26684, Z => n27443);
   U984 : BUF_X1 port map( A => n27281, Z => n27276);
   U985 : BUF_X1 port map( A => n26695, Z => n27281);
   U986 : BUF_X1 port map( A => n27371, Z => n27366);
   U987 : BUF_X1 port map( A => n26664, Z => n27371);
   U988 : BUF_X1 port map( A => n27365, Z => n27360);
   U989 : BUF_X1 port map( A => n26665, Z => n27365);
   U990 : BUF_X1 port map( A => n27359, Z => n27354);
   U991 : BUF_X1 port map( A => n26666, Z => n27359);
   U992 : BUF_X1 port map( A => n27353, Z => n27348);
   U993 : BUF_X1 port map( A => n26667, Z => n27353);
   U994 : BUF_X1 port map( A => n27347, Z => n27342);
   U995 : BUF_X1 port map( A => n26668, Z => n27347);
   U996 : BUF_X1 port map( A => n27341, Z => n27336);
   U997 : BUF_X1 port map( A => n26669, Z => n27341);
   U998 : BUF_X1 port map( A => n27335, Z => n27330);
   U999 : BUF_X1 port map( A => n26670, Z => n27335);
   U1000 : BUF_X1 port map( A => n27329, Z => n27324);
   U1001 : BUF_X1 port map( A => n26671, Z => n27329);
   U1002 : BUF_X1 port map( A => n27323, Z => n27318);
   U1003 : BUF_X1 port map( A => n26672, Z => n27323);
   U1004 : BUF_X1 port map( A => n27317, Z => n27312);
   U1005 : BUF_X1 port map( A => n26673, Z => n27317);
   U1006 : BUF_X1 port map( A => n27311, Z => n27306);
   U1007 : BUF_X1 port map( A => n26674, Z => n27311);
   U1008 : BUF_X1 port map( A => n27305, Z => n27300);
   U1009 : BUF_X1 port map( A => n26675, Z => n27305);
   U1010 : BUF_X1 port map( A => n27299, Z => n27294);
   U1011 : BUF_X1 port map( A => n26676, Z => n27299);
   U1012 : BUF_X1 port map( A => n27293, Z => n27288);
   U1013 : BUF_X1 port map( A => n26677, Z => n27293);
   U1014 : BUF_X1 port map( A => n27287, Z => n27282);
   U1015 : BUF_X1 port map( A => n26678, Z => n27287);
   U1016 : BUF_X1 port map( A => n27437, Z => n27432);
   U1017 : BUF_X1 port map( A => n26685, Z => n27437);
   U1018 : BUF_X1 port map( A => n27431, Z => n27426);
   U1019 : BUF_X1 port map( A => n26686, Z => n27431);
   U1020 : BUF_X1 port map( A => n27425, Z => n27420);
   U1021 : BUF_X1 port map( A => n26687, Z => n27425);
   U1022 : BUF_X1 port map( A => n27419, Z => n27414);
   U1023 : BUF_X1 port map( A => n26688, Z => n27419);
   U1024 : BUF_X1 port map( A => n27413, Z => n27408);
   U1025 : BUF_X1 port map( A => n26689, Z => n27413);
   U1026 : BUF_X1 port map( A => n27407, Z => n27402);
   U1027 : BUF_X1 port map( A => n26690, Z => n27407);
   U1028 : BUF_X1 port map( A => n27401, Z => n27396);
   U1029 : BUF_X1 port map( A => n26691, Z => n27401);
   U1030 : BUF_X1 port map( A => n27395, Z => n27390);
   U1031 : BUF_X1 port map( A => n26692, Z => n27395);
   U1032 : BUF_X1 port map( A => n27389, Z => n27384);
   U1033 : BUF_X1 port map( A => n26693, Z => n27389);
   U1034 : BUF_X1 port map( A => n27383, Z => n27378);
   U1035 : BUF_X1 port map( A => n26694, Z => n27383);
   U1036 : BUF_X1 port map( A => n27377, Z => n27372);
   U1037 : BUF_X1 port map( A => n26679, Z => n27377);
   U1038 : NOR3_X1 port map( A1 => add_rd2(0), A2 => add_rd2(1), A3 => n27713, 
                           ZN => n1235);
   U1039 : NOR3_X1 port map( A1 => n27704, A2 => add_rd2(2), A3 => n27712, ZN 
                           => n1236);
   U1040 : NOR3_X1 port map( A1 => add_rd2(1), A2 => add_rd2(2), A3 => n27704, 
                           ZN => n1243);
   U1041 : NOR2_X1 port map( A1 => add_rd1(3), A2 => add_rd1(4), ZN => n1854);
   U1042 : NOR2_X1 port map( A1 => n27718, A2 => add_rd1(4), ZN => n1853);
   U1043 : NOR3_X1 port map( A1 => add_rd1(1), A2 => add_rd1(2), A3 => 
                           add_rd1(0), ZN => n1861);
   U1044 : NOR3_X1 port map( A1 => add_rd1(0), A2 => add_rd1(1), A3 => n27717, 
                           ZN => n1855);
   U1045 : NOR2_X1 port map( A1 => n27719, A2 => add_rd1(3), ZN => n1872);
   U1046 : NOR3_X1 port map( A1 => add_rd2(0), A2 => add_rd2(2), A3 => n27712, 
                           ZN => n1234);
   U1047 : NOR3_X1 port map( A1 => add_rd1(1), A2 => add_rd1(2), A3 => n27715, 
                           ZN => n1864);
   U1048 : NOR3_X1 port map( A1 => add_rd2(1), A2 => add_rd2(2), A3 => 
                           add_rd2(0), ZN => n1238);
   U1049 : NOR3_X1 port map( A1 => n27712, A2 => add_rd2(0), A3 => n27713, ZN 
                           => n1233);
   U1050 : NOR3_X1 port map( A1 => add_rd1(0), A2 => add_rd1(2), A3 => n27716, 
                           ZN => n1858);
   U1051 : NOR3_X1 port map( A1 => n27716, A2 => add_rd1(0), A3 => n27717, ZN 
                           => n1857);
   U1052 : NOR3_X1 port map( A1 => n27715, A2 => add_rd1(2), A3 => n27716, ZN 
                           => n1852);
   U1053 : NOR3_X1 port map( A1 => n27715, A2 => add_rd1(1), A3 => n27717, ZN 
                           => n1860);
   U1054 : NOR3_X1 port map( A1 => n27704, A2 => add_rd2(1), A3 => n27713, ZN 
                           => n1239);
   U1055 : OAI221_X1 port map( B1 => n2547, B2 => n795_port, C1 => n2548, C2 =>
                           n796_port, A => n1125, ZN => n1120);
   U1056 : AOI22_X1 port map( A1 => n27707, A2 => n26696, B1 => n2546, B2 => 
                           n27701, ZN => n1125);
   U1057 : OAI221_X1 port map( B1 => n2551_port, B2 => n795_port, C1 => n2552, 
                           C2 => n796_port, A => n1107, ZN => n1102);
   U1058 : AOI22_X1 port map( A1 => n27707, A2 => n26697, B1 => n2550, B2 => 
                           n27701, ZN => n1107);
   U1059 : OAI221_X1 port map( B1 => n2555, B2 => n795_port, C1 => n2556, C2 =>
                           n796_port, A => n1089, ZN => n1084);
   U1060 : AOI22_X1 port map( A1 => n2553, A2 => n27707, B1 => n2554, B2 => 
                           n27701, ZN => n1089);
   U1061 : OAI221_X1 port map( B1 => n2559, B2 => n795_port, C1 => n2560, C2 =>
                           n796_port, A => n1071, ZN => n1066);
   U1062 : AOI22_X1 port map( A1 => n2557, A2 => n27707, B1 => n2558, B2 => 
                           n27701, ZN => n1071);
   U1063 : OAI221_X1 port map( B1 => n2563, B2 => n795_port, C1 => n2564, C2 =>
                           n796_port, A => n1053, ZN => n1048);
   U1064 : AOI22_X1 port map( A1 => n2561, A2 => n27707, B1 => n2562, B2 => 
                           n27701, ZN => n1053);
   U1065 : OAI221_X1 port map( B1 => n2567, B2 => n795_port, C1 => n2568, C2 =>
                           n796_port, A => n1017_port, ZN => n1012_port);
   U1066 : AOI22_X1 port map( A1 => n2565, A2 => n27707, B1 => n2566, B2 => 
                           n27701, ZN => n1017_port);
   U1067 : OAI221_X1 port map( B1 => n2571, B2 => n795_port, C1 => n2572, C2 =>
                           n796_port, A => n999_port, ZN => n994_port);
   U1068 : AOI22_X1 port map( A1 => n2569, A2 => n27707, B1 => n2570, B2 => 
                           n27701, ZN => n999_port);
   U1069 : OAI221_X1 port map( B1 => n2575, B2 => n795_port, C1 => n2576, C2 =>
                           n796_port, A => n981_port, ZN => n976_port);
   U1070 : AOI22_X1 port map( A1 => n2573, A2 => n27707, B1 => n2574, B2 => 
                           n27701, ZN => n981_port);
   U1071 : OAI221_X1 port map( B1 => n2579, B2 => n795_port, C1 => n2580, C2 =>
                           n796_port, A => n963_port, ZN => n958_port);
   U1072 : AOI22_X1 port map( A1 => n2577, A2 => n27707, B1 => n2578, B2 => 
                           n27701, ZN => n963_port);
   U1073 : OAI221_X1 port map( B1 => n2583_port, B2 => n795_port, C1 => n2584, 
                           C2 => n796_port, A => n945_port, ZN => n940_port);
   U1074 : AOI22_X1 port map( A1 => n2581, A2 => n27707, B1 => n2582, B2 => 
                           n27701, ZN => n945_port);
   U1075 : OAI221_X1 port map( B1 => n2587, B2 => n795_port, C1 => n2588, C2 =>
                           n796_port, A => n927_port, ZN => n922_port);
   U1076 : AOI22_X1 port map( A1 => n2585, A2 => n27707, B1 => n2586, B2 => 
                           n27701, ZN => n927_port);
   U1077 : OAI221_X1 port map( B1 => n2591, B2 => n795_port, C1 => n2592, C2 =>
                           n796_port, A => n909_port, ZN => n904_port);
   U1078 : AOI22_X1 port map( A1 => n2589, A2 => n27707, B1 => n2590, B2 => 
                           n27701, ZN => n909_port);
   U1079 : OAI221_X1 port map( B1 => n2595, B2 => n795_port, C1 => n2596, C2 =>
                           n796_port, A => n891_port, ZN => n886_port);
   U1080 : AOI22_X1 port map( A1 => n2593, A2 => n27707, B1 => n2594, B2 => 
                           n27701, ZN => n891_port);
   U1081 : OAI221_X1 port map( B1 => n2599, B2 => n795_port, C1 => n2600, C2 =>
                           n796_port, A => n873_port, ZN => n868_port);
   U1082 : AOI22_X1 port map( A1 => n2597, A2 => n27707, B1 => n2598, B2 => 
                           n27701, ZN => n873_port);
   U1083 : OAI221_X1 port map( B1 => n2603, B2 => n795_port, C1 => n2604, C2 =>
                           n796_port, A => n855_port, ZN => n850_port);
   U1084 : AOI22_X1 port map( A1 => n2601, A2 => n27707, B1 => n2602, B2 => 
                           n27701, ZN => n855_port);
   U1085 : OAI221_X1 port map( B1 => n2607, B2 => n795_port, C1 => n2608, C2 =>
                           n796_port, A => n819_port, ZN => n814_port);
   U1086 : AOI22_X1 port map( A1 => n2605, A2 => n27707, B1 => n2606, B2 => 
                           n27701, ZN => n819_port);
   U1087 : OAI221_X1 port map( B1 => n2611, B2 => n795_port, C1 => n2612, C2 =>
                           n796_port, A => n797_port, ZN => n790_port);
   U1088 : AOI22_X1 port map( A1 => n2609, A2 => n27707, B1 => n2610, B2 => 
                           n27701, ZN => n797_port);
   U1089 : OAI221_X1 port map( B1 => n25500, B2 => n651_port, C1 => n25259, C2 
                           => n652_port, A => n1242, ZN => n1228);
   U1090 : AOI22_X1 port map( A1 => n25434, A2 => n27703, B1 => n25179, B2 => 
                           n27702, ZN => n1242);
   U1091 : OAI221_X1 port map( B1 => n25501, B2 => n651_port, C1 => n25260, C2 
                           => n652_port, A => n1035_port, ZN => n1030_port);
   U1092 : AOI22_X1 port map( A1 => n25435, A2 => n27703, B1 => n25180, B2 => 
                           n27702, ZN => n1035_port);
   U1093 : OAI221_X1 port map( B1 => n25502, B2 => n651_port, C1 => n25261, C2 
                           => n652_port, A => n837_port, ZN => n832_port);
   U1094 : AOI22_X1 port map( A1 => n25436, A2 => n27703, B1 => n25181, B2 => 
                           n27702, ZN => n837_port);
   U1095 : OAI221_X1 port map( B1 => n25503, B2 => n651_port, C1 => n25262, C2 
                           => n652_port, A => n777_port, ZN => n772_port);
   U1096 : AOI22_X1 port map( A1 => n25437, A2 => n27703, B1 => n25182, B2 => 
                           n27702, ZN => n777_port);
   U1097 : OAI221_X1 port map( B1 => n25504, B2 => n651_port, C1 => n25263, C2 
                           => n652_port, A => n759_port, ZN => n754_port);
   U1098 : AOI22_X1 port map( A1 => n25438, A2 => n27703, B1 => n25183, B2 => 
                           n27702, ZN => n759_port);
   U1099 : OAI221_X1 port map( B1 => n25505, B2 => n651_port, C1 => n25264, C2 
                           => n652_port, A => n741_port, ZN => n736_port);
   U1100 : AOI22_X1 port map( A1 => n25439, A2 => n27703, B1 => n25184, B2 => 
                           n27702, ZN => n741_port);
   U1101 : OAI221_X1 port map( B1 => n25506, B2 => n651_port, C1 => n25265, C2 
                           => n652_port, A => n723_port, ZN => n718_port);
   U1102 : AOI22_X1 port map( A1 => n25440, A2 => n27703, B1 => n25185, B2 => 
                           n27702, ZN => n723_port);
   U1103 : OAI221_X1 port map( B1 => n25507, B2 => n651_port, C1 => n25266, C2 
                           => n652_port, A => n705_port, ZN => n700_port);
   U1104 : AOI22_X1 port map( A1 => n25441, A2 => n27703, B1 => n25186, B2 => 
                           n27702, ZN => n705_port);
   U1105 : OAI221_X1 port map( B1 => n25508, B2 => n651_port, C1 => n25267, C2 
                           => n652_port, A => n687_port, ZN => n682_port);
   U1106 : AOI22_X1 port map( A1 => n25442, A2 => n27703, B1 => n27702, B2 => 
                           n26593, ZN => n687_port);
   U1107 : OAI221_X1 port map( B1 => n25509, B2 => n651_port, C1 => n25268, C2 
                           => n652_port, A => n653_port, ZN => n638_port);
   U1108 : AOI22_X1 port map( A1 => n25443, A2 => n27703, B1 => n27702, B2 => 
                           n26594, ZN => n653_port);
   U1109 : OAI221_X1 port map( B1 => n25510, B2 => n651_port, C1 => n25269, C2 
                           => n652_port, A => n1215, ZN => n1210);
   U1110 : AOI22_X1 port map( A1 => n25444, A2 => n27703, B1 => n27702, B2 => 
                           n26595, ZN => n1215);
   U1111 : OAI221_X1 port map( B1 => n2142, B2 => n805_port, C1 => n2141, C2 =>
                           n806_port, A => n1025_port, ZN => n1020_port);
   U1112 : AOI22_X1 port map( A1 => n2139, A2 => n27708, B1 => n2140, B2 => 
                           n27709, ZN => n1025_port);
   U1113 : OAI221_X1 port map( B1 => n2149, B2 => n805_port, C1 => n2148, C2 =>
                           n806_port, A => n1007_port, ZN => n1002_port);
   U1114 : AOI22_X1 port map( A1 => n2146, A2 => n27708, B1 => n2147, B2 => 
                           n27709, ZN => n1007_port);
   U1115 : OAI221_X1 port map( B1 => n2156, B2 => n805_port, C1 => n2155, C2 =>
                           n806_port, A => n989_port, ZN => n984_port);
   U1116 : AOI22_X1 port map( A1 => n2153, A2 => n27708, B1 => n2154, B2 => 
                           n27709, ZN => n989_port);
   U1117 : OAI221_X1 port map( B1 => n2163, B2 => n805_port, C1 => n2162, C2 =>
                           n806_port, A => n971_port, ZN => n966_port);
   U1118 : AOI22_X1 port map( A1 => n2160, A2 => n27708, B1 => n2161, B2 => 
                           n27709, ZN => n971_port);
   U1119 : OAI221_X1 port map( B1 => n2170, B2 => n805_port, C1 => n2169, C2 =>
                           n806_port, A => n953_port, ZN => n948_port);
   U1120 : AOI22_X1 port map( A1 => n2167, A2 => n27708, B1 => n2168, B2 => 
                           n27709, ZN => n953_port);
   U1121 : OAI221_X1 port map( B1 => n2177, B2 => n805_port, C1 => n2176, C2 =>
                           n806_port, A => n935_port, ZN => n930_port);
   U1122 : AOI22_X1 port map( A1 => n2174, A2 => n27708, B1 => n2175, B2 => 
                           n27709, ZN => n935_port);
   U1123 : OAI221_X1 port map( B1 => n2184, B2 => n805_port, C1 => n2183, C2 =>
                           n806_port, A => n917_port, ZN => n912_port);
   U1124 : AOI22_X1 port map( A1 => n2181, A2 => n27708, B1 => n2182, B2 => 
                           n27709, ZN => n917_port);
   U1125 : OAI221_X1 port map( B1 => n2191, B2 => n805_port, C1 => n2190, C2 =>
                           n806_port, A => n899_port, ZN => n894_port);
   U1126 : AOI22_X1 port map( A1 => n2188, A2 => n27708, B1 => n2189, B2 => 
                           n27709, ZN => n899_port);
   U1127 : OAI221_X1 port map( B1 => n2198, B2 => n805_port, C1 => n2197, C2 =>
                           n806_port, A => n881_port, ZN => n876_port);
   U1128 : AOI22_X1 port map( A1 => n2195, A2 => n27708, B1 => n2196, B2 => 
                           n27709, ZN => n881_port);
   U1129 : OAI221_X1 port map( B1 => n2205, B2 => n805_port, C1 => n2204, C2 =>
                           n806_port, A => n863_port, ZN => n858_port);
   U1130 : AOI22_X1 port map( A1 => n2202, A2 => n27708, B1 => n2203, B2 => 
                           n27709, ZN => n863_port);
   U1131 : OAI221_X1 port map( B1 => n2212, B2 => n805_port, C1 => n2211, C2 =>
                           n806_port, A => n827_port, ZN => n822_port);
   U1132 : AOI22_X1 port map( A1 => n2209, A2 => n27708, B1 => n2210, B2 => 
                           n27709, ZN => n827_port);
   U1133 : OAI221_X1 port map( B1 => n2219, B2 => n805_port, C1 => n2218, C2 =>
                           n806_port, A => n807_port, ZN => n800_port);
   U1134 : AOI22_X1 port map( A1 => n2216, A2 => n27708, B1 => n2217, B2 => 
                           n27709, ZN => n807_port);
   U1135 : OAI221_X1 port map( B1 => n25250, B2 => n808_port, C1 => n25557, C2 
                           => n809_port, A => n972_port, ZN => n965_port);
   U1136 : AOI22_X1 port map( A1 => n25491, A2 => n27195, B1 => n25236, B2 => 
                           n27192, ZN => n972_port);
   U1137 : OAI221_X1 port map( B1 => n25251, B2 => n808_port, C1 => n25558, C2 
                           => n809_port, A => n954_port, ZN => n947_port);
   U1138 : AOI22_X1 port map( A1 => n25492, A2 => n27195, B1 => n25237, B2 => 
                           n27192, ZN => n954_port);
   U1139 : OAI221_X1 port map( B1 => n25252, B2 => n808_port, C1 => n25559, C2 
                           => n809_port, A => n936_port, ZN => n929_port);
   U1140 : AOI22_X1 port map( A1 => n25493, A2 => n27195, B1 => n25238, B2 => 
                           n27192, ZN => n936_port);
   U1141 : OAI221_X1 port map( B1 => n25253, B2 => n808_port, C1 => n25560, C2 
                           => n809_port, A => n918_port, ZN => n911_port);
   U1142 : AOI22_X1 port map( A1 => n25494, A2 => n27195, B1 => n25239, B2 => 
                           n27192, ZN => n918_port);
   U1143 : OAI221_X1 port map( B1 => n25254, B2 => n808_port, C1 => n25561, C2 
                           => n809_port, A => n900_port, ZN => n893_port);
   U1144 : AOI22_X1 port map( A1 => n25495, A2 => n27195, B1 => n25240, B2 => 
                           n27192, ZN => n900_port);
   U1145 : OAI221_X1 port map( B1 => n25255, B2 => n808_port, C1 => n25562, C2 
                           => n809_port, A => n882_port, ZN => n875_port);
   U1146 : AOI22_X1 port map( A1 => n25496, A2 => n27195, B1 => n25241, B2 => 
                           n27192, ZN => n882_port);
   U1147 : OAI221_X1 port map( B1 => n25256, B2 => n808_port, C1 => n25563, C2 
                           => n809_port, A => n864_port, ZN => n857_port);
   U1148 : AOI22_X1 port map( A1 => n25497, A2 => n27195, B1 => n25242, B2 => 
                           n27192, ZN => n864_port);
   U1149 : OAI221_X1 port map( B1 => n25257, B2 => n808_port, C1 => n25564, C2 
                           => n809_port, A => n828_port, ZN => n821_port);
   U1150 : AOI22_X1 port map( A1 => n25498, A2 => n27195, B1 => n25243, B2 => 
                           n27192, ZN => n828_port);
   U1151 : OAI221_X1 port map( B1 => n25258, B2 => n808_port, C1 => n25565, C2 
                           => n809_port, A => n810_port, ZN => n799_port);
   U1152 : AOI22_X1 port map( A1 => n25499, A2 => n27195, B1 => n25244, B2 => 
                           n27192, ZN => n810_port);
   U1153 : OAI221_X1 port map( B1 => n2359_port, B2 => n27273, C1 => n2360, C2 
                           => n27269, A => n1231, ZN => n1230);
   U1154 : AOI22_X1 port map( A1 => n2423_port, A2 => n27265, B1 => n2424, B2 
                           => n27261, ZN => n1231);
   U1155 : OAI221_X1 port map( B1 => n27225, B2 => n26600, C1 => n27221, C2 => 
                           n26327, A => n1249, ZN => n1248);
   U1156 : AOI22_X1 port map( A1 => regs_13_0_port, A2 => n27217, B1 => 
                           regs_5_0_port, B2 => n27213, ZN => n1249);
   U1157 : OAI221_X1 port map( B1 => n2361, B2 => n27274, C1 => n2362, C2 => 
                           n27270, A => n1033_port, ZN => n1032_port);
   U1158 : AOI22_X1 port map( A1 => n2425, A2 => n27265, B1 => n2426, B2 => 
                           n27261, ZN => n1033_port);
   U1159 : OAI221_X1 port map( B1 => n27225, B2 => n26601, C1 => n27222, C2 => 
                           n26328, A => n1041_port, ZN => n1040_port);
   U1160 : AOI22_X1 port map( A1 => regs_13_1_port, A2 => n27217, B1 => 
                           regs_5_1_port, B2 => n27213, ZN => n1041_port);
   U1161 : OAI221_X1 port map( B1 => n2363, B2 => n27275, C1 => n2364, C2 => 
                           n27271, A => n835_port, ZN => n834_port);
   U1162 : AOI22_X1 port map( A1 => n2427, A2 => n27266, B1 => n2428, B2 => 
                           n27262, ZN => n835_port);
   U1163 : OAI221_X1 port map( B1 => n27226, B2 => n26602, C1 => n27223, C2 => 
                           n26329, A => n843_port, ZN => n842_port);
   U1164 : AOI22_X1 port map( A1 => regs_13_2_port, A2 => n27218, B1 => 
                           regs_5_2_port, B2 => n27214, ZN => n843_port);
   U1165 : OAI221_X1 port map( B1 => n2365, B2 => n27275, C1 => n2366, C2 => 
                           n27271, A => n775_port, ZN => n774_port);
   U1166 : AOI22_X1 port map( A1 => n2429, A2 => n27267, B1 => n2430, B2 => 
                           n27263, ZN => n775_port);
   U1167 : OAI221_X1 port map( B1 => n27227, B2 => n26603, C1 => n27223, C2 => 
                           n26330, A => n783_port, ZN => n782_port);
   U1168 : AOI22_X1 port map( A1 => regs_13_3_port, A2 => n27219, B1 => 
                           regs_5_3_port, B2 => n27215, ZN => n783_port);
   U1169 : OAI221_X1 port map( B1 => n2367, B2 => n27275, C1 => n2368, C2 => 
                           n27271, A => n757_port, ZN => n756_port);
   U1170 : AOI22_X1 port map( A1 => n2431, A2 => n27267, B1 => n2432, B2 => 
                           n27263, ZN => n757_port);
   U1171 : OAI221_X1 port map( B1 => n27227, B2 => n26604, C1 => n27223, C2 => 
                           n26331, A => n765_port, ZN => n764_port);
   U1172 : AOI22_X1 port map( A1 => regs_13_4_port, A2 => n27219, B1 => 
                           regs_5_4_port, B2 => n27215, ZN => n765_port);
   U1173 : OAI221_X1 port map( B1 => n2369, B2 => n27275, C1 => n2370, C2 => 
                           n27271, A => n739_port, ZN => n738_port);
   U1174 : AOI22_X1 port map( A1 => n2433, A2 => n27267, B1 => n2434, B2 => 
                           n27263, ZN => n739_port);
   U1175 : OAI221_X1 port map( B1 => n27227, B2 => n26605, C1 => n27223, C2 => 
                           n26332, A => n747_port, ZN => n746_port);
   U1176 : AOI22_X1 port map( A1 => regs_13_5_port, A2 => n27219, B1 => 
                           regs_5_5_port, B2 => n27215, ZN => n747_port);
   U1177 : OAI221_X1 port map( B1 => n2371, B2 => n27275, C1 => n2372, C2 => 
                           n27271, A => n721_port, ZN => n720_port);
   U1178 : AOI22_X1 port map( A1 => n2435, A2 => n27267, B1 => n2436, B2 => 
                           n27263, ZN => n721_port);
   U1179 : OAI221_X1 port map( B1 => n27227, B2 => n26606, C1 => n27223, C2 => 
                           n26333, A => n729_port, ZN => n728_port);
   U1180 : AOI22_X1 port map( A1 => regs_13_6_port, A2 => n27219, B1 => 
                           regs_5_6_port, B2 => n27215, ZN => n729_port);
   U1181 : OAI221_X1 port map( B1 => n2373, B2 => n27275, C1 => n2374, C2 => 
                           n27271, A => n703_port, ZN => n702_port);
   U1182 : AOI22_X1 port map( A1 => n2437, A2 => n27267, B1 => n2438, B2 => 
                           n27263, ZN => n703_port);
   U1183 : OAI221_X1 port map( B1 => n27227, B2 => n26607, C1 => n27223, C2 => 
                           n26334, A => n711_port, ZN => n710_port);
   U1184 : AOI22_X1 port map( A1 => regs_13_7_port, A2 => n27219, B1 => 
                           regs_5_7_port, B2 => n27215, ZN => n711_port);
   U1185 : OAI221_X1 port map( B1 => n2375, B2 => n27275, C1 => n2376, C2 => 
                           n27271, A => n685_port, ZN => n684_port);
   U1186 : AOI22_X1 port map( A1 => n2439, A2 => n27267, B1 => n2440, B2 => 
                           n27263, ZN => n685_port);
   U1187 : OAI221_X1 port map( B1 => n27227, B2 => n26608, C1 => n27223, C2 => 
                           n26335, A => n693_port, ZN => n692_port);
   U1188 : AOI22_X1 port map( A1 => regs_13_8_port, A2 => n27219, B1 => 
                           regs_5_8_port, B2 => n27215, ZN => n693_port);
   U1189 : OAI221_X1 port map( B1 => n2377, B2 => n27275, C1 => n2378, C2 => 
                           n27271, A => n643_port, ZN => n640_port);
   U1190 : AOI22_X1 port map( A1 => n2441, A2 => n27267, B1 => n2442, B2 => 
                           n27263, ZN => n643_port);
   U1191 : OAI221_X1 port map( B1 => n27227, B2 => n26609, C1 => n27223, C2 => 
                           n26336, A => n665_port, ZN => n662_port);
   U1192 : AOI22_X1 port map( A1 => regs_13_9_port, A2 => n27219, B1 => 
                           regs_5_9_port, B2 => n27215, ZN => n665_port);
   U1193 : OAI221_X1 port map( B1 => n2379, B2 => n27273, C1 => n2380, C2 => 
                           n27269, A => n1213, ZN => n1212);
   U1194 : AOI22_X1 port map( A1 => n2443, A2 => n27265, B1 => n2444, B2 => 
                           n27261, ZN => n1213);
   U1195 : OAI221_X1 port map( B1 => n27225, B2 => n26610, C1 => n27221, C2 => 
                           n26337, A => n1221, ZN => n1220);
   U1196 : AOI22_X1 port map( A1 => regs_13_10_port, A2 => n27217, B1 => 
                           regs_5_10_port, B2 => n27213, ZN => n1221);
   U1197 : OAI221_X1 port map( B1 => n2381, B2 => n27273, C1 => n2382, C2 => 
                           n27269, A => n1194, ZN => n1193);
   U1198 : AOI22_X1 port map( A1 => n2445, A2 => n27265, B1 => n2446, B2 => 
                           n27261, ZN => n1194);
   U1199 : OAI221_X1 port map( B1 => n27225, B2 => n26611, C1 => n27221, C2 => 
                           n26338, A => n1203, ZN => n1202);
   U1200 : AOI22_X1 port map( A1 => regs_13_11_port, A2 => n27217, B1 => 
                           regs_5_11_port, B2 => n27213, ZN => n1203);
   U1201 : OAI221_X1 port map( B1 => n2383, B2 => n27273, C1 => n2384, C2 => 
                           n27269, A => n1176, ZN => n1175);
   U1202 : AOI22_X1 port map( A1 => n2447, A2 => n27265, B1 => n2448, B2 => 
                           n27261, ZN => n1176);
   U1203 : OAI221_X1 port map( B1 => n27225, B2 => n26612, C1 => n27221, C2 => 
                           n26339, A => n1185, ZN => n1184);
   U1204 : AOI22_X1 port map( A1 => regs_13_12_port, A2 => n27217, B1 => 
                           regs_5_12_port, B2 => n27213, ZN => n1185);
   U1205 : OAI221_X1 port map( B1 => n2385, B2 => n27273, C1 => n2386, C2 => 
                           n27269, A => n1158, ZN => n1157);
   U1206 : AOI22_X1 port map( A1 => n2449, A2 => n27265, B1 => n2450, B2 => 
                           n27261, ZN => n1158);
   U1207 : OAI221_X1 port map( B1 => n27225, B2 => n26613, C1 => n27221, C2 => 
                           n26340, A => n1167, ZN => n1166);
   U1208 : AOI22_X1 port map( A1 => regs_13_13_port, A2 => n27217, B1 => 
                           regs_5_13_port, B2 => n27213, ZN => n1167);
   U1209 : OAI221_X1 port map( B1 => n2387, B2 => n27273, C1 => n2388, C2 => 
                           n27269, A => n1140, ZN => n1139);
   U1210 : AOI22_X1 port map( A1 => n2451, A2 => n27265, B1 => n2452, B2 => 
                           n27261, ZN => n1140);
   U1211 : OAI221_X1 port map( B1 => n27225, B2 => n26614, C1 => n27221, C2 => 
                           n26341, A => n1149, ZN => n1148);
   U1212 : AOI22_X1 port map( A1 => regs_13_14_port, A2 => n27217, B1 => 
                           regs_5_14_port, B2 => n27213, ZN => n1149);
   U1213 : OAI221_X1 port map( B1 => n2389, B2 => n27273, C1 => n2390, C2 => 
                           n27269, A => n1123, ZN => n1122);
   U1214 : AOI22_X1 port map( A1 => n2453, A2 => n27265, B1 => n2454, B2 => 
                           n27261, ZN => n1123);
   U1215 : OAI221_X1 port map( B1 => n27225, B2 => n26615, C1 => n27221, C2 => 
                           n26342, A => n1131, ZN => n1130);
   U1216 : AOI22_X1 port map( A1 => regs_13_15_port, A2 => n27217, B1 => 
                           regs_5_15_port, B2 => n27213, ZN => n1131);
   U1217 : OAI221_X1 port map( B1 => n2391_port, B2 => n27273, C1 => n2392, C2 
                           => n27269, A => n1105, ZN => n1104);
   U1218 : AOI22_X1 port map( A1 => n2455_port, A2 => n27265, B1 => n2456, B2 
                           => n27261, ZN => n1105);
   U1219 : OAI221_X1 port map( B1 => n27225, B2 => n26616, C1 => n27221, C2 => 
                           n26343, A => n1113, ZN => n1112);
   U1220 : AOI22_X1 port map( A1 => regs_13_16_port, A2 => n27217, B1 => 
                           regs_5_16_port, B2 => n27213, ZN => n1113);
   U1221 : OAI221_X1 port map( B1 => n2393, B2 => n27273, C1 => n2394, C2 => 
                           n27269, A => n1087, ZN => n1086);
   U1222 : AOI22_X1 port map( A1 => n2457, A2 => n27265, B1 => n2458, B2 => 
                           n27261, ZN => n1087);
   U1223 : OAI221_X1 port map( B1 => n27225, B2 => n26617, C1 => n27221, C2 => 
                           n26344, A => n1095, ZN => n1094);
   U1224 : AOI22_X1 port map( A1 => regs_13_17_port, A2 => n27217, B1 => 
                           regs_5_17_port, B2 => n27213, ZN => n1095);
   U1225 : OAI221_X1 port map( B1 => n2395, B2 => n27273, C1 => n2396, C2 => 
                           n27269, A => n1069, ZN => n1068);
   U1226 : AOI22_X1 port map( A1 => n2459, A2 => n27265, B1 => n2460, B2 => 
                           n27261, ZN => n1069);
   U1227 : OAI221_X1 port map( B1 => n27225, B2 => n26618, C1 => n27221, C2 => 
                           n26345, A => n1077, ZN => n1076);
   U1228 : AOI22_X1 port map( A1 => regs_13_18_port, A2 => n27217, B1 => 
                           regs_5_18_port, B2 => n27213, ZN => n1077);
   U1229 : OAI221_X1 port map( B1 => n2397, B2 => n27273, C1 => n2398, C2 => 
                           n27269, A => n1051, ZN => n1050);
   U1230 : AOI22_X1 port map( A1 => n2461, A2 => n27265, B1 => n2462, B2 => 
                           n27261, ZN => n1051);
   U1231 : OAI221_X1 port map( B1 => n27225, B2 => n26619, C1 => n27221, C2 => 
                           n26346, A => n1059, ZN => n1058);
   U1232 : AOI22_X1 port map( A1 => regs_13_19_port, A2 => n27217, B1 => 
                           regs_5_19_port, B2 => n27213, ZN => n1059);
   U1233 : OAI221_X1 port map( B1 => n2399, B2 => n27274, C1 => n2400, C2 => 
                           n27270, A => n1015_port, ZN => n1014_port);
   U1234 : AOI22_X1 port map( A1 => n2463, A2 => n27266, B1 => n2464, B2 => 
                           n27262, ZN => n1015_port);
   U1235 : OAI221_X1 port map( B1 => n27226, B2 => n26620, C1 => n27222, C2 => 
                           n26347, A => n1023_port, ZN => n1022_port);
   U1236 : AOI22_X1 port map( A1 => regs_13_20_port, A2 => n27218, B1 => 
                           regs_5_20_port, B2 => n27214, ZN => n1023_port);
   U1237 : OAI221_X1 port map( B1 => n2401, B2 => n27274, C1 => n2402, C2 => 
                           n27270, A => n997_port, ZN => n996_port);
   U1238 : AOI22_X1 port map( A1 => n2465, A2 => n27266, B1 => n2466, B2 => 
                           n27262, ZN => n997_port);
   U1239 : OAI221_X1 port map( B1 => n27226, B2 => n26621, C1 => n27222, C2 => 
                           n26348, A => n1005_port, ZN => n1004_port);
   U1240 : AOI22_X1 port map( A1 => regs_13_21_port, A2 => n27218, B1 => 
                           regs_5_21_port, B2 => n27214, ZN => n1005_port);
   U1241 : OAI221_X1 port map( B1 => n2403, B2 => n27274, C1 => n2404, C2 => 
                           n27270, A => n979_port, ZN => n978_port);
   U1242 : AOI22_X1 port map( A1 => n2467, A2 => n27266, B1 => n2468, B2 => 
                           n27262, ZN => n979_port);
   U1243 : OAI221_X1 port map( B1 => n27226, B2 => n26622, C1 => n27222, C2 => 
                           n26349, A => n987_port, ZN => n986_port);
   U1244 : AOI22_X1 port map( A1 => regs_13_22_port, A2 => n27218, B1 => 
                           regs_5_22_port, B2 => n27214, ZN => n987_port);
   U1245 : OAI221_X1 port map( B1 => n2405, B2 => n27274, C1 => n2406, C2 => 
                           n27270, A => n961_port, ZN => n960_port);
   U1246 : AOI22_X1 port map( A1 => n2469, A2 => n27266, B1 => n2470, B2 => 
                           n27262, ZN => n961_port);
   U1247 : OAI221_X1 port map( B1 => n27226, B2 => n26623, C1 => n27222, C2 => 
                           n26350, A => n969_port, ZN => n968_port);
   U1248 : AOI22_X1 port map( A1 => regs_13_23_port, A2 => n27218, B1 => 
                           regs_5_23_port, B2 => n27214, ZN => n969_port);
   U1249 : OAI221_X1 port map( B1 => n2407, B2 => n27274, C1 => n2408, C2 => 
                           n27270, A => n943_port, ZN => n942_port);
   U1250 : AOI22_X1 port map( A1 => n2471, A2 => n27266, B1 => n2472, B2 => 
                           n27262, ZN => n943_port);
   U1251 : OAI221_X1 port map( B1 => n27226, B2 => n26624, C1 => n27222, C2 => 
                           n26351, A => n951_port, ZN => n950_port);
   U1252 : AOI22_X1 port map( A1 => regs_13_24_port, A2 => n27218, B1 => 
                           regs_5_24_port, B2 => n27214, ZN => n951_port);
   U1253 : OAI221_X1 port map( B1 => n2409, B2 => n27274, C1 => n2410, C2 => 
                           n27270, A => n925_port, ZN => n924_port);
   U1254 : AOI22_X1 port map( A1 => n2473, A2 => n27266, B1 => n2474, B2 => 
                           n27262, ZN => n925_port);
   U1255 : OAI221_X1 port map( B1 => n27226, B2 => n26625, C1 => n27222, C2 => 
                           n26352, A => n933_port, ZN => n932_port);
   U1256 : AOI22_X1 port map( A1 => regs_13_25_port, A2 => n27218, B1 => 
                           regs_5_25_port, B2 => n27214, ZN => n933_port);
   U1257 : OAI221_X1 port map( B1 => n2411, B2 => n27274, C1 => n2412, C2 => 
                           n27270, A => n907_port, ZN => n906_port);
   U1258 : AOI22_X1 port map( A1 => n2475, A2 => n27266, B1 => n2476, B2 => 
                           n27262, ZN => n907_port);
   U1259 : OAI221_X1 port map( B1 => n27226, B2 => n26626, C1 => n27222, C2 => 
                           n26353, A => n915_port, ZN => n914_port);
   U1260 : AOI22_X1 port map( A1 => regs_13_26_port, A2 => n27218, B1 => 
                           regs_5_26_port, B2 => n27214, ZN => n915_port);
   U1261 : OAI221_X1 port map( B1 => n2413, B2 => n27274, C1 => n2414, C2 => 
                           n27270, A => n889_port, ZN => n888_port);
   U1262 : AOI22_X1 port map( A1 => n2477, A2 => n27266, B1 => n2478, B2 => 
                           n27262, ZN => n889_port);
   U1263 : OAI221_X1 port map( B1 => n27226, B2 => n26627, C1 => n27222, C2 => 
                           n26354, A => n897_port, ZN => n896_port);
   U1264 : AOI22_X1 port map( A1 => regs_13_27_port, A2 => n27218, B1 => 
                           regs_5_27_port, B2 => n27214, ZN => n897_port);
   U1265 : OAI221_X1 port map( B1 => n2415, B2 => n27274, C1 => n2416, C2 => 
                           n27270, A => n871_port, ZN => n870_port);
   U1266 : AOI22_X1 port map( A1 => n2479, A2 => n27266, B1 => n2480, B2 => 
                           n27262, ZN => n871_port);
   U1267 : OAI221_X1 port map( B1 => n27226, B2 => n26628, C1 => n27222, C2 => 
                           n26355, A => n879_port, ZN => n878_port);
   U1268 : AOI22_X1 port map( A1 => regs_13_28_port, A2 => n27218, B1 => 
                           regs_5_28_port, B2 => n27214, ZN => n879_port);
   U1269 : OAI221_X1 port map( B1 => n2417, B2 => n27274, C1 => n2418, C2 => 
                           n27270, A => n853_port, ZN => n852_port);
   U1270 : AOI22_X1 port map( A1 => n2481, A2 => n27266, B1 => n2482, B2 => 
                           n27262, ZN => n853_port);
   U1271 : OAI221_X1 port map( B1 => n27226, B2 => n26629, C1 => n27222, C2 => 
                           n26356, A => n861_port, ZN => n860_port);
   U1272 : AOI22_X1 port map( A1 => regs_13_29_port, A2 => n27218, B1 => 
                           regs_5_29_port, B2 => n27214, ZN => n861_port);
   U1273 : OAI221_X1 port map( B1 => n2419, B2 => n27275, C1 => n2420, C2 => 
                           n27271, A => n817_port, ZN => n816_port);
   U1274 : AOI22_X1 port map( A1 => n2483, A2 => n27266, B1 => n2484, B2 => 
                           n27262, ZN => n817_port);
   U1275 : OAI221_X1 port map( B1 => n27226, B2 => n26630, C1 => n27223, C2 => 
                           n26357, A => n825_port, ZN => n824_port);
   U1276 : AOI22_X1 port map( A1 => regs_13_30_port, A2 => n27218, B1 => 
                           regs_5_30_port, B2 => n27214, ZN => n825_port);
   U1277 : OAI221_X1 port map( B1 => n2421, B2 => n27275, C1 => n2422, C2 => 
                           n27271, A => n793_port, ZN => n792_port);
   U1278 : AOI22_X1 port map( A1 => n2485, A2 => n27267, B1 => n2486, B2 => 
                           n27263, ZN => n793_port);
   U1279 : OAI221_X1 port map( B1 => n27227, B2 => n26631, C1 => n27223, C2 => 
                           n26358, A => n803_port, ZN => n802_port);
   U1280 : AOI22_X1 port map( A1 => regs_13_31_port, A2 => n27219, B1 => 
                           regs_5_31_port, B2 => n27215, ZN => n803_port);
   U1281 : OAI221_X1 port map( B1 => n26475, B2 => n27187, C1 => n26907, C2 => 
                           n27183, A => n1851, ZN => n1850);
   U1282 : AOI22_X1 port map( A1 => n27179, A2 => n26391, B1 => n27175, B2 => 
                           n26730, ZN => n1851);
   U1283 : OAI221_X1 port map( B1 => n2359_port, B2 => n27123, C1 => n2360, C2 
                           => n27119, A => n1869, ZN => n1868);
   U1284 : AOI22_X1 port map( A1 => n27115, A2 => n2423_port, B1 => n27111, B2 
                           => n2424, ZN => n1869);
   U1285 : OAI221_X1 port map( B1 => n26476, B2 => n27188, C1 => n26908, C2 => 
                           n27184, A => n1653, ZN => n1652);
   U1286 : AOI22_X1 port map( A1 => n27180, A2 => n26392, B1 => n27176, B2 => 
                           n26731, ZN => n1653);
   U1287 : OAI221_X1 port map( B1 => n2361, B2 => n27124, C1 => n2362, C2 => 
                           n27120, A => n1661, ZN => n1660);
   U1288 : AOI22_X1 port map( A1 => n27116, A2 => n2425, B1 => n27112, B2 => 
                           n2426, ZN => n1661);
   U1289 : OAI221_X1 port map( B1 => n26477, B2 => n27189, C1 => n26909, C2 => 
                           n27185, A => n1455, ZN => n1454);
   U1290 : AOI22_X1 port map( A1 => n27181, A2 => n26393, B1 => n27177, B2 => 
                           n26732, ZN => n1455);
   U1291 : OAI221_X1 port map( B1 => n2363, B2 => n27125, C1 => n2364, C2 => 
                           n27121, A => n1463, ZN => n1462);
   U1292 : AOI22_X1 port map( A1 => n27117, A2 => n2427, B1 => n27113, B2 => 
                           n2428, ZN => n1463);
   U1293 : OAI221_X1 port map( B1 => n26478, B2 => n27189, C1 => n26910, C2 => 
                           n27185, A => n1401, ZN => n1400);
   U1294 : AOI22_X1 port map( A1 => n27181, A2 => n26394, B1 => n27177, B2 => 
                           n26733, ZN => n1401);
   U1295 : OAI221_X1 port map( B1 => n2365, B2 => n27125, C1 => n2366, C2 => 
                           n27121, A => n1409, ZN => n1408);
   U1296 : AOI22_X1 port map( A1 => n27117, A2 => n2429, B1 => n27113, B2 => 
                           n2430, ZN => n1409);
   U1297 : OAI221_X1 port map( B1 => n26479, B2 => n27189, C1 => n26911, C2 => 
                           n27185, A => n1383, ZN => n1382);
   U1298 : AOI22_X1 port map( A1 => n27181, A2 => n26395, B1 => n27177, B2 => 
                           n26734, ZN => n1383);
   U1299 : OAI221_X1 port map( B1 => n2367, B2 => n27125, C1 => n2368, C2 => 
                           n27121, A => n1391, ZN => n1390);
   U1300 : AOI22_X1 port map( A1 => n27117, A2 => n2431, B1 => n27113, B2 => 
                           n2432, ZN => n1391);
   U1301 : OAI221_X1 port map( B1 => n26480, B2 => n27189, C1 => n26912, C2 => 
                           n27185, A => n1365, ZN => n1364);
   U1302 : AOI22_X1 port map( A1 => n27181, A2 => n26396, B1 => n27177, B2 => 
                           n26735, ZN => n1365);
   U1303 : OAI221_X1 port map( B1 => n2369, B2 => n27125, C1 => n2370, C2 => 
                           n27121, A => n1373, ZN => n1372);
   U1304 : AOI22_X1 port map( A1 => n27117, A2 => n2433, B1 => n27113, B2 => 
                           n2434, ZN => n1373);
   U1305 : OAI221_X1 port map( B1 => n26481, B2 => n27189, C1 => n26913, C2 => 
                           n27185, A => n1347, ZN => n1346);
   U1306 : AOI22_X1 port map( A1 => n27181, A2 => n26397, B1 => n27177, B2 => 
                           n26736, ZN => n1347);
   U1307 : OAI221_X1 port map( B1 => n2371, B2 => n27125, C1 => n2372, C2 => 
                           n27121, A => n1355, ZN => n1354);
   U1308 : AOI22_X1 port map( A1 => n27117, A2 => n2435, B1 => n27113, B2 => 
                           n2436, ZN => n1355);
   U1309 : OAI221_X1 port map( B1 => n26482, B2 => n27189, C1 => n26914, C2 => 
                           n27185, A => n1329, ZN => n1328);
   U1310 : AOI22_X1 port map( A1 => n27181, A2 => n26398, B1 => n27177, B2 => 
                           n26737, ZN => n1329);
   U1311 : OAI221_X1 port map( B1 => n2373, B2 => n27125, C1 => n2374, C2 => 
                           n27121, A => n1337, ZN => n1336);
   U1312 : AOI22_X1 port map( A1 => n27117, A2 => n2437, B1 => n27113, B2 => 
                           n2438, ZN => n1337);
   U1313 : OAI221_X1 port map( B1 => n26483, B2 => n27189, C1 => n26915, C2 => 
                           n27185, A => n1311, ZN => n1310);
   U1314 : AOI22_X1 port map( A1 => n27181, A2 => n26399, B1 => n27177, B2 => 
                           n26738, ZN => n1311);
   U1315 : OAI221_X1 port map( B1 => n2375, B2 => n27125, C1 => n2376, C2 => 
                           n27121, A => n1319, ZN => n1318);
   U1316 : AOI22_X1 port map( A1 => n27117, A2 => n2439, B1 => n27113, B2 => 
                           n2440, ZN => n1319);
   U1317 : OAI221_X1 port map( B1 => n26484, B2 => n27189, C1 => n26916, C2 => 
                           n27185, A => n1263, ZN => n1260);
   U1318 : AOI22_X1 port map( A1 => n27181, A2 => n26400, B1 => n27177, B2 => 
                           n26739, ZN => n1263);
   U1319 : OAI221_X1 port map( B1 => n2377, B2 => n27125, C1 => n2378, C2 => 
                           n27121, A => n1287, ZN => n1284);
   U1320 : AOI22_X1 port map( A1 => n27117, A2 => n2441, B1 => n27113, B2 => 
                           n2442, ZN => n1287);
   U1321 : OAI221_X1 port map( B1 => n26485, B2 => n27187, C1 => n26917, C2 => 
                           n27183, A => n1833, ZN => n1832);
   U1322 : AOI22_X1 port map( A1 => n27179, A2 => n26401, B1 => n27175, B2 => 
                           n26740, ZN => n1833);
   U1323 : OAI221_X1 port map( B1 => n2379, B2 => n27123, C1 => n2380, C2 => 
                           n27119, A => n1841, ZN => n1840);
   U1324 : AOI22_X1 port map( A1 => n27115, A2 => n2443, B1 => n27111, B2 => 
                           n2444, ZN => n1841);
   U1325 : OAI221_X1 port map( B1 => n26486, B2 => n27187, C1 => n26918, C2 => 
                           n27183, A => n1815, ZN => n1814);
   U1326 : AOI22_X1 port map( A1 => n27179, A2 => n26402, B1 => n27175, B2 => 
                           n26741, ZN => n1815);
   U1327 : OAI221_X1 port map( B1 => n2381, B2 => n27123, C1 => n2382, C2 => 
                           n27119, A => n1823, ZN => n1822);
   U1328 : AOI22_X1 port map( A1 => n27115, A2 => n2445, B1 => n27111, B2 => 
                           n2446, ZN => n1823);
   U1329 : OAI221_X1 port map( B1 => n26487, B2 => n27187, C1 => n26919, C2 => 
                           n27183, A => n1797, ZN => n1796);
   U1330 : AOI22_X1 port map( A1 => n27179, A2 => n26403, B1 => n27175, B2 => 
                           n26742, ZN => n1797);
   U1331 : OAI221_X1 port map( B1 => n2383, B2 => n27123, C1 => n2384, C2 => 
                           n27119, A => n1805, ZN => n1804);
   U1332 : AOI22_X1 port map( A1 => n27115, A2 => n2447, B1 => n27111, B2 => 
                           n2448, ZN => n1805);
   U1333 : OAI221_X1 port map( B1 => n26488, B2 => n27187, C1 => n26920, C2 => 
                           n27183, A => n1779, ZN => n1778);
   U1334 : AOI22_X1 port map( A1 => n27179, A2 => n26404, B1 => n27175, B2 => 
                           n26743, ZN => n1779);
   U1335 : OAI221_X1 port map( B1 => n2385, B2 => n27123, C1 => n2386, C2 => 
                           n27119, A => n1787, ZN => n1786);
   U1336 : AOI22_X1 port map( A1 => n27115, A2 => n2449, B1 => n27111, B2 => 
                           n2450, ZN => n1787);
   U1337 : OAI221_X1 port map( B1 => n26489, B2 => n27187, C1 => n26921, C2 => 
                           n27183, A => n1761, ZN => n1760);
   U1338 : AOI22_X1 port map( A1 => n27179, A2 => n26405, B1 => n27175, B2 => 
                           n26744, ZN => n1761);
   U1339 : OAI221_X1 port map( B1 => n2387, B2 => n27123, C1 => n2388, C2 => 
                           n27119, A => n1769, ZN => n1768);
   U1340 : AOI22_X1 port map( A1 => n27115, A2 => n2451, B1 => n27111, B2 => 
                           n2452, ZN => n1769);
   U1341 : OAI221_X1 port map( B1 => n26490, B2 => n27187, C1 => n26922, C2 => 
                           n27183, A => n1743, ZN => n1742);
   U1342 : AOI22_X1 port map( A1 => n27179, A2 => n26406, B1 => n27175, B2 => 
                           n26745, ZN => n1743);
   U1343 : OAI221_X1 port map( B1 => n2389, B2 => n27123, C1 => n2390, C2 => 
                           n27119, A => n1751, ZN => n1750);
   U1344 : AOI22_X1 port map( A1 => n27115, A2 => n2453, B1 => n27111, B2 => 
                           n2454, ZN => n1751);
   U1345 : OAI221_X1 port map( B1 => n26491, B2 => n27187, C1 => n26923, C2 => 
                           n27183, A => n1725, ZN => n1724);
   U1346 : AOI22_X1 port map( A1 => n27179, A2 => n26407, B1 => n27175, B2 => 
                           n26746, ZN => n1725);
   U1347 : OAI221_X1 port map( B1 => n2391_port, B2 => n27123, C1 => n2392, C2 
                           => n27119, A => n1733, ZN => n1732);
   U1348 : AOI22_X1 port map( A1 => n27115, A2 => n2455_port, B1 => n27111, B2 
                           => n2456, ZN => n1733);
   U1349 : OAI221_X1 port map( B1 => n26492, B2 => n27187, C1 => n26924, C2 => 
                           n27183, A => n1707, ZN => n1706);
   U1350 : AOI22_X1 port map( A1 => n27179, A2 => n26408, B1 => n27175, B2 => 
                           n26747, ZN => n1707);
   U1351 : OAI221_X1 port map( B1 => n2393, B2 => n27123, C1 => n2394, C2 => 
                           n27119, A => n1715, ZN => n1714);
   U1352 : AOI22_X1 port map( A1 => n27115, A2 => n2457, B1 => n27111, B2 => 
                           n2458, ZN => n1715);
   U1353 : OAI221_X1 port map( B1 => n26493, B2 => n27187, C1 => n26925, C2 => 
                           n27183, A => n1689, ZN => n1688);
   U1354 : AOI22_X1 port map( A1 => n27179, A2 => n26409, B1 => n27175, B2 => 
                           n26748, ZN => n1689);
   U1355 : OAI221_X1 port map( B1 => n2395, B2 => n27123, C1 => n2396, C2 => 
                           n27119, A => n1697, ZN => n1696);
   U1356 : AOI22_X1 port map( A1 => n27115, A2 => n2459, B1 => n27111, B2 => 
                           n2460, ZN => n1697);
   U1357 : OAI221_X1 port map( B1 => n26494, B2 => n27187, C1 => n26926, C2 => 
                           n27183, A => n1671, ZN => n1670);
   U1358 : AOI22_X1 port map( A1 => n27179, A2 => n26410, B1 => n27175, B2 => 
                           n26749, ZN => n1671);
   U1359 : OAI221_X1 port map( B1 => n2397, B2 => n27123, C1 => n2398, C2 => 
                           n27119, A => n1679, ZN => n1678);
   U1360 : AOI22_X1 port map( A1 => n27115, A2 => n2461, B1 => n27111, B2 => 
                           n2462, ZN => n1679);
   U1361 : OAI221_X1 port map( B1 => n26495, B2 => n27188, C1 => n26927, C2 => 
                           n27184, A => n1635, ZN => n1634);
   U1362 : AOI22_X1 port map( A1 => n27180, A2 => n26411, B1 => n27176, B2 => 
                           n26750, ZN => n1635);
   U1363 : OAI221_X1 port map( B1 => n2399, B2 => n27124, C1 => n2400, C2 => 
                           n27120, A => n1643, ZN => n1642);
   U1364 : AOI22_X1 port map( A1 => n27116, A2 => n2463, B1 => n27112, B2 => 
                           n2464, ZN => n1643);
   U1365 : OAI221_X1 port map( B1 => n26496, B2 => n27188, C1 => n26928, C2 => 
                           n27184, A => n1617, ZN => n1616);
   U1366 : AOI22_X1 port map( A1 => n27180, A2 => n26412, B1 => n27176, B2 => 
                           n26751, ZN => n1617);
   U1367 : OAI221_X1 port map( B1 => n2401, B2 => n27124, C1 => n2402, C2 => 
                           n27120, A => n1625, ZN => n1624);
   U1368 : AOI22_X1 port map( A1 => n27116, A2 => n2465, B1 => n27112, B2 => 
                           n2466, ZN => n1625);
   U1369 : OAI221_X1 port map( B1 => n26497, B2 => n27188, C1 => n26929, C2 => 
                           n27184, A => n1599, ZN => n1598);
   U1370 : AOI22_X1 port map( A1 => n27180, A2 => n26413, B1 => n27176, B2 => 
                           n26752, ZN => n1599);
   U1371 : OAI221_X1 port map( B1 => n2403, B2 => n27124, C1 => n2404, C2 => 
                           n27120, A => n1607, ZN => n1606);
   U1372 : AOI22_X1 port map( A1 => n27116, A2 => n2467, B1 => n27112, B2 => 
                           n2468, ZN => n1607);
   U1373 : OAI221_X1 port map( B1 => n25557, B2 => n27188, C1 => n25250, C2 => 
                           n27184, A => n1581, ZN => n1580);
   U1374 : AOI22_X1 port map( A1 => n27180, A2 => n25491, B1 => n27176, B2 => 
                           n25236, ZN => n1581);
   U1375 : OAI221_X1 port map( B1 => n2405, B2 => n27124, C1 => n2406, C2 => 
                           n27120, A => n1589, ZN => n1588);
   U1376 : AOI22_X1 port map( A1 => n27116, A2 => n2469, B1 => n27112, B2 => 
                           n2470, ZN => n1589);
   U1377 : OAI221_X1 port map( B1 => n25558, B2 => n27188, C1 => n25251, C2 => 
                           n27184, A => n1563, ZN => n1562);
   U1378 : AOI22_X1 port map( A1 => n27180, A2 => n25492, B1 => n27176, B2 => 
                           n25237, ZN => n1563);
   U1379 : OAI221_X1 port map( B1 => n2407, B2 => n27124, C1 => n2408, C2 => 
                           n27120, A => n1571, ZN => n1570);
   U1380 : AOI22_X1 port map( A1 => n27116, A2 => n2471, B1 => n27112, B2 => 
                           n2472, ZN => n1571);
   U1381 : OAI221_X1 port map( B1 => n25559, B2 => n27188, C1 => n25252, C2 => 
                           n27184, A => n1545, ZN => n1544);
   U1382 : AOI22_X1 port map( A1 => n27180, A2 => n25493, B1 => n27176, B2 => 
                           n25238, ZN => n1545);
   U1383 : OAI221_X1 port map( B1 => n2409, B2 => n27124, C1 => n2410, C2 => 
                           n27120, A => n1553, ZN => n1552);
   U1384 : AOI22_X1 port map( A1 => n27116, A2 => n2473, B1 => n27112, B2 => 
                           n2474, ZN => n1553);
   U1385 : OAI221_X1 port map( B1 => n25560, B2 => n27188, C1 => n25253, C2 => 
                           n27184, A => n1527, ZN => n1526);
   U1386 : AOI22_X1 port map( A1 => n27180, A2 => n25494, B1 => n27176, B2 => 
                           n25239, ZN => n1527);
   U1387 : OAI221_X1 port map( B1 => n2411, B2 => n27124, C1 => n2412, C2 => 
                           n27120, A => n1535, ZN => n1534);
   U1388 : AOI22_X1 port map( A1 => n27116, A2 => n2475, B1 => n27112, B2 => 
                           n2476, ZN => n1535);
   U1389 : OAI221_X1 port map( B1 => n25561, B2 => n27188, C1 => n25254, C2 => 
                           n27184, A => n1509, ZN => n1508);
   U1390 : AOI22_X1 port map( A1 => n27180, A2 => n25495, B1 => n27176, B2 => 
                           n25240, ZN => n1509);
   U1391 : OAI221_X1 port map( B1 => n2413, B2 => n27124, C1 => n2414, C2 => 
                           n27120, A => n1517, ZN => n1516);
   U1392 : AOI22_X1 port map( A1 => n27116, A2 => n2477, B1 => n27112, B2 => 
                           n2478, ZN => n1517);
   U1393 : OAI221_X1 port map( B1 => n25562, B2 => n27188, C1 => n25255, C2 => 
                           n27184, A => n1491, ZN => n1490);
   U1394 : AOI22_X1 port map( A1 => n27180, A2 => n25496, B1 => n27176, B2 => 
                           n25241, ZN => n1491);
   U1395 : OAI221_X1 port map( B1 => n2415, B2 => n27124, C1 => n2416, C2 => 
                           n27120, A => n1499, ZN => n1498);
   U1396 : AOI22_X1 port map( A1 => n27116, A2 => n2479, B1 => n27112, B2 => 
                           n2480, ZN => n1499);
   U1397 : OAI221_X1 port map( B1 => n25563, B2 => n27188, C1 => n25256, C2 => 
                           n27184, A => n1473, ZN => n1472);
   U1398 : AOI22_X1 port map( A1 => n27180, A2 => n25497, B1 => n27176, B2 => 
                           n25242, ZN => n1473);
   U1399 : OAI221_X1 port map( B1 => n2417, B2 => n27124, C1 => n2418, C2 => 
                           n27120, A => n1481, ZN => n1480);
   U1400 : AOI22_X1 port map( A1 => n27116, A2 => n2481, B1 => n27112, B2 => 
                           n2482, ZN => n1481);
   U1401 : OAI221_X1 port map( B1 => n25564, B2 => n27189, C1 => n25257, C2 => 
                           n27185, A => n1437, ZN => n1436);
   U1402 : AOI22_X1 port map( A1 => n27181, A2 => n25498, B1 => n27177, B2 => 
                           n25243, ZN => n1437);
   U1403 : OAI221_X1 port map( B1 => n2419, B2 => n27125, C1 => n2420, C2 => 
                           n27121, A => n1445, ZN => n1444);
   U1404 : AOI22_X1 port map( A1 => n27117, A2 => n2483, B1 => n27113, B2 => 
                           n2484, ZN => n1445);
   U1405 : OAI221_X1 port map( B1 => n25565, B2 => n27189, C1 => n25258, C2 => 
                           n27185, A => n1419, ZN => n1418);
   U1406 : AOI22_X1 port map( A1 => n27181, A2 => n25499, B1 => n27177, B2 => 
                           n25244, ZN => n1419);
   U1407 : OAI221_X1 port map( B1 => n2421, B2 => n27125, C1 => n2422, C2 => 
                           n27121, A => n1427, ZN => n1426);
   U1408 : AOI22_X1 port map( A1 => n27117, A2 => n2485, B1 => n27113, B2 => 
                           n2486, ZN => n1427);
   U1409 : OAI221_X1 port map( B1 => n25532, B2 => n27171, C1 => n25291, C2 => 
                           n27167, A => n1856, ZN => n1849);
   U1410 : AOI22_X1 port map( A1 => n27163, A2 => n25466, B1 => n27159, B2 => 
                           n25211, ZN => n1856);
   U1411 : OAI221_X1 port map( B1 => n25533, B2 => n27172, C1 => n25292, C2 => 
                           n27168, A => n1654, ZN => n1651);
   U1412 : AOI22_X1 port map( A1 => n27164, A2 => n25467, B1 => n27160, B2 => 
                           n25212, ZN => n1654);
   U1413 : OAI221_X1 port map( B1 => n25534, B2 => n27173, C1 => n25293, C2 => 
                           n27169, A => n1456, ZN => n1453);
   U1414 : AOI22_X1 port map( A1 => n27165, A2 => n25468, B1 => n27161, B2 => 
                           n25213, ZN => n1456);
   U1415 : OAI221_X1 port map( B1 => n25535, B2 => n27173, C1 => n25294, C2 => 
                           n27169, A => n1402, ZN => n1399);
   U1416 : AOI22_X1 port map( A1 => n27165, A2 => n25469, B1 => n27161, B2 => 
                           n25214, ZN => n1402);
   U1417 : OAI221_X1 port map( B1 => n25536, B2 => n27173, C1 => n25295, C2 => 
                           n27169, A => n1384, ZN => n1381);
   U1418 : AOI22_X1 port map( A1 => n27165, A2 => n25470, B1 => n27161, B2 => 
                           n25215, ZN => n1384);
   U1419 : OAI221_X1 port map( B1 => n25537, B2 => n27173, C1 => n25296, C2 => 
                           n27169, A => n1366, ZN => n1363);
   U1420 : AOI22_X1 port map( A1 => n27165, A2 => n25471, B1 => n27161, B2 => 
                           n25216, ZN => n1366);
   U1421 : OAI221_X1 port map( B1 => n25538, B2 => n27173, C1 => n25297, C2 => 
                           n27169, A => n1348, ZN => n1345);
   U1422 : AOI22_X1 port map( A1 => n27165, A2 => n25472, B1 => n27161, B2 => 
                           n25217, ZN => n1348);
   U1423 : OAI221_X1 port map( B1 => n25539, B2 => n27173, C1 => n25298, C2 => 
                           n27169, A => n1330, ZN => n1327);
   U1424 : AOI22_X1 port map( A1 => n27165, A2 => n25473, B1 => n27161, B2 => 
                           n25218, ZN => n1330);
   U1425 : OAI221_X1 port map( B1 => n25540, B2 => n27173, C1 => n25299, C2 => 
                           n27169, A => n1312, ZN => n1309);
   U1426 : AOI22_X1 port map( A1 => n27165, A2 => n25474, B1 => n27161, B2 => 
                           n25219, ZN => n1312);
   U1427 : OAI221_X1 port map( B1 => n25541, B2 => n27173, C1 => n25300, C2 => 
                           n27169, A => n1268, ZN => n1259);
   U1428 : AOI22_X1 port map( A1 => n27165, A2 => n25475, B1 => n27161, B2 => 
                           n25220, ZN => n1268);
   U1429 : OAI221_X1 port map( B1 => n25542, B2 => n27171, C1 => n25301, C2 => 
                           n27167, A => n1834, ZN => n1831);
   U1430 : AOI22_X1 port map( A1 => n27163, A2 => n25476, B1 => n27159, B2 => 
                           n25221, ZN => n1834);
   U1431 : OAI221_X1 port map( B1 => n25543, B2 => n27171, C1 => n25302, C2 => 
                           n27167, A => n1816, ZN => n1813);
   U1432 : AOI22_X1 port map( A1 => n27163, A2 => n25477, B1 => n27159, B2 => 
                           n25222, ZN => n1816);
   U1433 : OAI221_X1 port map( B1 => n25544, B2 => n27171, C1 => n25303, C2 => 
                           n27167, A => n1798, ZN => n1795);
   U1434 : AOI22_X1 port map( A1 => n27163, A2 => n25478, B1 => n27159, B2 => 
                           n25223, ZN => n1798);
   U1435 : OAI221_X1 port map( B1 => n25545, B2 => n27171, C1 => n25304, C2 => 
                           n27167, A => n1780, ZN => n1777);
   U1436 : AOI22_X1 port map( A1 => n27163, A2 => n25479, B1 => n27159, B2 => 
                           n25224, ZN => n1780);
   U1437 : OAI221_X1 port map( B1 => n25546, B2 => n27171, C1 => n25305, C2 => 
                           n27167, A => n1762, ZN => n1759);
   U1438 : AOI22_X1 port map( A1 => n27163, A2 => n25480, B1 => n27159, B2 => 
                           n25225, ZN => n1762);
   U1439 : OAI221_X1 port map( B1 => n25547, B2 => n27171, C1 => n25306, C2 => 
                           n27167, A => n1744, ZN => n1741);
   U1440 : AOI22_X1 port map( A1 => n27163, A2 => n25481, B1 => n27159, B2 => 
                           n25226, ZN => n1744);
   U1441 : OAI221_X1 port map( B1 => n25548, B2 => n27171, C1 => n25307, C2 => 
                           n27167, A => n1726, ZN => n1723);
   U1442 : AOI22_X1 port map( A1 => n27163, A2 => n25482, B1 => n27159, B2 => 
                           n25227, ZN => n1726);
   U1443 : OAI221_X1 port map( B1 => n25549, B2 => n27171, C1 => n25308, C2 => 
                           n27167, A => n1708, ZN => n1705);
   U1444 : AOI22_X1 port map( A1 => n27163, A2 => n25483, B1 => n27159, B2 => 
                           n25228, ZN => n1708);
   U1445 : OAI221_X1 port map( B1 => n25550, B2 => n27171, C1 => n25309, C2 => 
                           n27167, A => n1690, ZN => n1687);
   U1446 : AOI22_X1 port map( A1 => n27163, A2 => n25484, B1 => n27159, B2 => 
                           n25229, ZN => n1690);
   U1447 : OAI221_X1 port map( B1 => n25551, B2 => n27171, C1 => n25310, C2 => 
                           n27167, A => n1672, ZN => n1669);
   U1448 : AOI22_X1 port map( A1 => n27163, A2 => n25485, B1 => n27159, B2 => 
                           n25230, ZN => n1672);
   U1449 : OAI221_X1 port map( B1 => n2081, B2 => n27257, C1 => n27253, C2 => 
                           n26930, A => n1237, ZN => n1229);
   U1450 : AOI22_X1 port map( A1 => n2079, A2 => n27249, B1 => n2080, B2 => 
                           n27245, ZN => n1237);
   U1451 : OAI221_X1 port map( B1 => n27209, B2 => n26632, C1 => n27205, C2 => 
                           n26359, A => n1252, ZN => n1247);
   U1452 : AOI22_X1 port map( A1 => regs_15_0_port, A2 => n27201, B1 => 
                           regs_7_0_port, B2 => n27197, ZN => n1252);
   U1453 : OAI221_X1 port map( B1 => n2084, B2 => n27258, C1 => n27254, C2 => 
                           n26931, A => n1034_port, ZN => n1031_port);
   U1454 : AOI22_X1 port map( A1 => n2082, A2 => n27249, B1 => n2083, B2 => 
                           n27245, ZN => n1034_port);
   U1455 : OAI221_X1 port map( B1 => n27209, B2 => n26633, C1 => n27206, C2 => 
                           n26360, A => n1042_port, ZN => n1039_port);
   U1456 : AOI22_X1 port map( A1 => regs_15_1_port, A2 => n27201, B1 => 
                           regs_7_1_port, B2 => n27197, ZN => n1042_port);
   U1457 : OAI221_X1 port map( B1 => n2087, B2 => n27259, C1 => n27255, C2 => 
                           n26932, A => n836_port, ZN => n833_port);
   U1458 : AOI22_X1 port map( A1 => n2085, A2 => n27250, B1 => n2086, B2 => 
                           n27246, ZN => n836_port);
   U1459 : OAI221_X1 port map( B1 => n27210, B2 => n26634, C1 => n27207, C2 => 
                           n26361, A => n844_port, ZN => n841_port);
   U1460 : AOI22_X1 port map( A1 => regs_15_2_port, A2 => n27202, B1 => 
                           regs_7_2_port, B2 => n27198, ZN => n844_port);
   U1461 : OAI221_X1 port map( B1 => n2090, B2 => n27259, C1 => n27255, C2 => 
                           n26933, A => n776_port, ZN => n773_port);
   U1462 : AOI22_X1 port map( A1 => n2088, A2 => n27251, B1 => n2089, B2 => 
                           n27247, ZN => n776_port);
   U1463 : OAI221_X1 port map( B1 => n27211, B2 => n26635, C1 => n27207, C2 => 
                           n26362, A => n784_port, ZN => n781_port);
   U1464 : AOI22_X1 port map( A1 => regs_15_3_port, A2 => n27203, B1 => 
                           regs_7_3_port, B2 => n27199, ZN => n784_port);
   U1465 : OAI221_X1 port map( B1 => n2093, B2 => n27259, C1 => n27255, C2 => 
                           n26934, A => n758_port, ZN => n755_port);
   U1466 : AOI22_X1 port map( A1 => n2091, A2 => n27251, B1 => n2092, B2 => 
                           n27247, ZN => n758_port);
   U1467 : OAI221_X1 port map( B1 => n27211, B2 => n26636, C1 => n27207, C2 => 
                           n26363, A => n766_port, ZN => n763_port);
   U1468 : AOI22_X1 port map( A1 => regs_15_4_port, A2 => n27203, B1 => 
                           regs_7_4_port, B2 => n27199, ZN => n766_port);
   U1469 : OAI221_X1 port map( B1 => n2096, B2 => n27259, C1 => n27255, C2 => 
                           n26935, A => n740_port, ZN => n737_port);
   U1470 : AOI22_X1 port map( A1 => n2094, A2 => n27251, B1 => n2095, B2 => 
                           n27247, ZN => n740_port);
   U1471 : OAI221_X1 port map( B1 => n27211, B2 => n26637, C1 => n27207, C2 => 
                           n26364, A => n748_port, ZN => n745_port);
   U1472 : AOI22_X1 port map( A1 => regs_15_5_port, A2 => n27203, B1 => 
                           regs_7_5_port, B2 => n27199, ZN => n748_port);
   U1473 : OAI221_X1 port map( B1 => n2099, B2 => n27259, C1 => n27255, C2 => 
                           n26936, A => n722_port, ZN => n719_port);
   U1474 : AOI22_X1 port map( A1 => n2097, A2 => n27251, B1 => n2098, B2 => 
                           n27247, ZN => n722_port);
   U1475 : OAI221_X1 port map( B1 => n27211, B2 => n26638, C1 => n27207, C2 => 
                           n26365, A => n730_port, ZN => n727_port);
   U1476 : AOI22_X1 port map( A1 => regs_15_6_port, A2 => n27203, B1 => 
                           regs_7_6_port, B2 => n27199, ZN => n730_port);
   U1477 : OAI221_X1 port map( B1 => n2102, B2 => n27259, C1 => n27255, C2 => 
                           n26937, A => n704_port, ZN => n701_port);
   U1478 : AOI22_X1 port map( A1 => n2100, A2 => n27251, B1 => n2101, B2 => 
                           n27247, ZN => n704_port);
   U1479 : OAI221_X1 port map( B1 => n27211, B2 => n26639, C1 => n27207, C2 => 
                           n26366, A => n712_port, ZN => n709_port);
   U1480 : AOI22_X1 port map( A1 => regs_15_7_port, A2 => n27203, B1 => 
                           regs_7_7_port, B2 => n27199, ZN => n712_port);
   U1481 : OAI221_X1 port map( B1 => n2105, B2 => n27259, C1 => n27255, C2 => 
                           n26938, A => n686_port, ZN => n683_port);
   U1482 : AOI22_X1 port map( A1 => n2103, A2 => n27251, B1 => n2104, B2 => 
                           n27247, ZN => n686_port);
   U1483 : OAI221_X1 port map( B1 => n27211, B2 => n26640, C1 => n27207, C2 => 
                           n26367, A => n694_port, ZN => n691_port);
   U1484 : AOI22_X1 port map( A1 => regs_15_8_port, A2 => n27203, B1 => 
                           regs_7_8_port, B2 => n27199, ZN => n694_port);
   U1485 : OAI221_X1 port map( B1 => n2108, B2 => n27259, C1 => n27255, C2 => 
                           n26939, A => n648_port, ZN => n639_port);
   U1486 : AOI22_X1 port map( A1 => n2106, A2 => n27251, B1 => n2107, B2 => 
                           n27247, ZN => n648_port);
   U1487 : OAI221_X1 port map( B1 => n27211, B2 => n26641, C1 => n27207, C2 => 
                           n26368, A => n670_port, ZN => n661_port);
   U1488 : AOI22_X1 port map( A1 => regs_15_9_port, A2 => n27203, B1 => 
                           regs_7_9_port, B2 => n27199, ZN => n670_port);
   U1489 : OAI221_X1 port map( B1 => n2111, B2 => n27257, C1 => n27253, C2 => 
                           n26940, A => n1214, ZN => n1211);
   U1490 : AOI22_X1 port map( A1 => n2109, A2 => n27249, B1 => n2110, B2 => 
                           n27245, ZN => n1214);
   U1491 : OAI221_X1 port map( B1 => n27209, B2 => n26642, C1 => n27205, C2 => 
                           n26369, A => n1222, ZN => n1219);
   U1492 : AOI22_X1 port map( A1 => regs_15_10_port, A2 => n27201, B1 => 
                           regs_7_10_port, B2 => n27197, ZN => n1222);
   U1493 : OAI221_X1 port map( B1 => n2114, B2 => n27257, C1 => n27253, C2 => 
                           n26941, A => n1195, ZN => n1192);
   U1494 : AOI22_X1 port map( A1 => n2112, A2 => n27249, B1 => n2113, B2 => 
                           n27245, ZN => n1195);
   U1495 : OAI221_X1 port map( B1 => n27209, B2 => n26643, C1 => n27205, C2 => 
                           n26370, A => n1204, ZN => n1201);
   U1496 : AOI22_X1 port map( A1 => regs_15_11_port, A2 => n27201, B1 => 
                           regs_7_11_port, B2 => n27197, ZN => n1204);
   U1497 : OAI221_X1 port map( B1 => n2117, B2 => n27257, C1 => n27253, C2 => 
                           n26942, A => n1177, ZN => n1174);
   U1498 : AOI22_X1 port map( A1 => n2115, A2 => n27249, B1 => n2116, B2 => 
                           n27245, ZN => n1177);
   U1499 : OAI221_X1 port map( B1 => n27209, B2 => n26644, C1 => n27205, C2 => 
                           n26371, A => n1186, ZN => n1183);
   U1500 : AOI22_X1 port map( A1 => regs_15_12_port, A2 => n27201, B1 => 
                           regs_7_12_port, B2 => n27197, ZN => n1186);
   U1501 : OAI221_X1 port map( B1 => n2120, B2 => n27257, C1 => n27253, C2 => 
                           n26943, A => n1159, ZN => n1156);
   U1502 : AOI22_X1 port map( A1 => n2118, A2 => n27249, B1 => n2119, B2 => 
                           n27245, ZN => n1159);
   U1503 : OAI221_X1 port map( B1 => n27209, B2 => n26645, C1 => n27205, C2 => 
                           n26372, A => n1168, ZN => n1165);
   U1504 : AOI22_X1 port map( A1 => regs_15_13_port, A2 => n27201, B1 => 
                           regs_7_13_port, B2 => n27197, ZN => n1168);
   U1505 : OAI221_X1 port map( B1 => n2123, B2 => n27257, C1 => n27253, C2 => 
                           n26944, A => n1141, ZN => n1138);
   U1506 : AOI22_X1 port map( A1 => n2121, A2 => n27249, B1 => n2122, B2 => 
                           n27245, ZN => n1141);
   U1507 : OAI221_X1 port map( B1 => n27209, B2 => n26646, C1 => n27205, C2 => 
                           n26373, A => n1150, ZN => n1147);
   U1508 : AOI22_X1 port map( A1 => regs_15_14_port, A2 => n27201, B1 => 
                           regs_7_14_port, B2 => n27197, ZN => n1150);
   U1509 : OAI221_X1 port map( B1 => n2126, B2 => n27257, C1 => n27253, C2 => 
                           n26945, A => n1124, ZN => n1121);
   U1510 : AOI22_X1 port map( A1 => n2124, A2 => n27249, B1 => n2125, B2 => 
                           n27245, ZN => n1124);
   U1511 : OAI221_X1 port map( B1 => n27209, B2 => n26647, C1 => n27205, C2 => 
                           n26374, A => n1132, ZN => n1129);
   U1512 : AOI22_X1 port map( A1 => regs_15_15_port, A2 => n27201, B1 => 
                           regs_7_15_port, B2 => n27197, ZN => n1132);
   U1513 : OAI221_X1 port map( B1 => n2129, B2 => n27257, C1 => n27253, C2 => 
                           n26946, A => n1106, ZN => n1103);
   U1514 : AOI22_X1 port map( A1 => n2127, A2 => n27249, B1 => n2128, B2 => 
                           n27245, ZN => n1106);
   U1515 : OAI221_X1 port map( B1 => n27209, B2 => n26648, C1 => n27205, C2 => 
                           n26375, A => n1114, ZN => n1111);
   U1516 : AOI22_X1 port map( A1 => regs_15_16_port, A2 => n27201, B1 => 
                           regs_7_16_port, B2 => n27197, ZN => n1114);
   U1517 : OAI221_X1 port map( B1 => n2132, B2 => n27257, C1 => n27253, C2 => 
                           n26947, A => n1088, ZN => n1085);
   U1518 : AOI22_X1 port map( A1 => n2130, A2 => n27249, B1 => n2131, B2 => 
                           n27245, ZN => n1088);
   U1519 : OAI221_X1 port map( B1 => n27209, B2 => n26649, C1 => n27205, C2 => 
                           n26376, A => n1096, ZN => n1093);
   U1520 : AOI22_X1 port map( A1 => regs_15_17_port, A2 => n27201, B1 => 
                           regs_7_17_port, B2 => n27197, ZN => n1096);
   U1521 : OAI221_X1 port map( B1 => n2135, B2 => n27257, C1 => n27253, C2 => 
                           n26948, A => n1070, ZN => n1067);
   U1522 : AOI22_X1 port map( A1 => n2133, A2 => n27249, B1 => n2134, B2 => 
                           n27245, ZN => n1070);
   U1523 : OAI221_X1 port map( B1 => n27209, B2 => n26650, C1 => n27205, C2 => 
                           n26377, A => n1078, ZN => n1075);
   U1524 : AOI22_X1 port map( A1 => regs_15_18_port, A2 => n27201, B1 => 
                           regs_7_18_port, B2 => n27197, ZN => n1078);
   U1525 : OAI221_X1 port map( B1 => n2138, B2 => n27257, C1 => n27253, C2 => 
                           n26949, A => n1052, ZN => n1049);
   U1526 : AOI22_X1 port map( A1 => n2136, A2 => n27249, B1 => n2137, B2 => 
                           n27245, ZN => n1052);
   U1527 : OAI221_X1 port map( B1 => n27209, B2 => n26651, C1 => n27205, C2 => 
                           n26378, A => n1060, ZN => n1057);
   U1528 : AOI22_X1 port map( A1 => regs_15_19_port, A2 => n27201, B1 => 
                           regs_7_19_port, B2 => n27197, ZN => n1060);
   U1529 : OAI221_X1 port map( B1 => n2145, B2 => n27258, C1 => n27254, C2 => 
                           n26950, A => n1016_port, ZN => n1013_port);
   U1530 : AOI22_X1 port map( A1 => n2143, A2 => n27250, B1 => n2144, B2 => 
                           n27246, ZN => n1016_port);
   U1531 : OAI221_X1 port map( B1 => n27210, B2 => n26652, C1 => n27206, C2 => 
                           n26379, A => n1024_port, ZN => n1021_port);
   U1532 : AOI22_X1 port map( A1 => regs_15_20_port, A2 => n27202, B1 => 
                           regs_7_20_port, B2 => n27198, ZN => n1024_port);
   U1533 : OAI221_X1 port map( B1 => n2152, B2 => n27258, C1 => n27254, C2 => 
                           n26951, A => n998_port, ZN => n995_port);
   U1534 : AOI22_X1 port map( A1 => n2150, A2 => n27250, B1 => n2151, B2 => 
                           n27246, ZN => n998_port);
   U1535 : OAI221_X1 port map( B1 => n27210, B2 => n26653, C1 => n27206, C2 => 
                           n26380, A => n1006_port, ZN => n1003_port);
   U1536 : AOI22_X1 port map( A1 => regs_15_21_port, A2 => n27202, B1 => 
                           regs_7_21_port, B2 => n27198, ZN => n1006_port);
   U1537 : OAI221_X1 port map( B1 => n2159, B2 => n27258, C1 => n27254, C2 => 
                           n26952, A => n980_port, ZN => n977_port);
   U1538 : AOI22_X1 port map( A1 => n2157, A2 => n27250, B1 => n2158, B2 => 
                           n27246, ZN => n980_port);
   U1539 : OAI221_X1 port map( B1 => n27210, B2 => n26654, C1 => n27206, C2 => 
                           n26381, A => n988_port, ZN => n985_port);
   U1540 : AOI22_X1 port map( A1 => regs_15_22_port, A2 => n27202, B1 => 
                           regs_7_22_port, B2 => n27198, ZN => n988_port);
   U1541 : OAI221_X1 port map( B1 => n2166_port, B2 => n27258, C1 => n27254, C2
                           => n26953, A => n962_port, ZN => n959_port);
   U1542 : AOI22_X1 port map( A1 => n2164, A2 => n27250, B1 => n2165, B2 => 
                           n27246, ZN => n962_port);
   U1543 : OAI221_X1 port map( B1 => n2173, B2 => n27258, C1 => n27254, C2 => 
                           n26954, A => n944_port, ZN => n941_port);
   U1544 : AOI22_X1 port map( A1 => n2171, A2 => n27250, B1 => n2172, B2 => 
                           n27246, ZN => n944_port);
   U1545 : OAI221_X1 port map( B1 => n2180, B2 => n27258, C1 => n27254, C2 => 
                           n26955, A => n926_port, ZN => n923_port);
   U1546 : AOI22_X1 port map( A1 => n2178, A2 => n27250, B1 => n2179, B2 => 
                           n27246, ZN => n926_port);
   U1547 : OAI221_X1 port map( B1 => n2187, B2 => n27258, C1 => n27254, C2 => 
                           n26956, A => n908_port, ZN => n905_port);
   U1548 : AOI22_X1 port map( A1 => n2185, A2 => n27250, B1 => n2186, B2 => 
                           n27246, ZN => n908_port);
   U1549 : OAI221_X1 port map( B1 => n2194, B2 => n27258, C1 => n27254, C2 => 
                           n26957, A => n890_port, ZN => n887_port);
   U1550 : AOI22_X1 port map( A1 => n2192, A2 => n27250, B1 => n2193, B2 => 
                           n27246, ZN => n890_port);
   U1551 : OAI221_X1 port map( B1 => n2201, B2 => n27258, C1 => n27254, C2 => 
                           n26958, A => n872_port, ZN => n869_port);
   U1552 : AOI22_X1 port map( A1 => n2199_port, A2 => n27250, B1 => n2200, B2 
                           => n27246, ZN => n872_port);
   U1553 : OAI221_X1 port map( B1 => n2208, B2 => n27258, C1 => n27254, C2 => 
                           n26959, A => n854_port, ZN => n851_port);
   U1554 : AOI22_X1 port map( A1 => n2206, A2 => n27250, B1 => n2207, B2 => 
                           n27246, ZN => n854_port);
   U1555 : OAI221_X1 port map( B1 => n2215, B2 => n27259, C1 => n27255, C2 => 
                           n26960, A => n818_port, ZN => n815_port);
   U1556 : AOI22_X1 port map( A1 => n2213, A2 => n27250, B1 => n2214, B2 => 
                           n27246, ZN => n818_port);
   U1557 : OAI221_X1 port map( B1 => n2222, B2 => n27259, C1 => n27255, C2 => 
                           n26961, A => n794_port, ZN => n791_port);
   U1558 : AOI22_X1 port map( A1 => n2220, A2 => n27251, B1 => n2221, B2 => 
                           n27247, ZN => n794_port);
   U1559 : OAI221_X1 port map( B1 => n26530, B2 => n27107, C1 => n26846, C2 => 
                           n27103, A => n1871, ZN => n1867);
   U1560 : AOI22_X1 port map( A1 => n27099, A2 => n26698, B1 => n27095, B2 => 
                           regs_18_0_port, ZN => n1871);
   U1561 : OAI221_X1 port map( B1 => n26531, B2 => n27108, C1 => n26847, C2 => 
                           n27104, A => n1662, ZN => n1659);
   U1562 : AOI22_X1 port map( A1 => n27100, A2 => n26699, B1 => n27096, B2 => 
                           regs_18_1_port, ZN => n1662);
   U1563 : OAI221_X1 port map( B1 => n26532, B2 => n27109, C1 => n26848, C2 => 
                           n27105, A => n1464, ZN => n1461);
   U1564 : AOI22_X1 port map( A1 => n27101, A2 => n26700, B1 => n27097, B2 => 
                           regs_18_2_port, ZN => n1464);
   U1565 : OAI221_X1 port map( B1 => n26533, B2 => n27109, C1 => n26849, C2 => 
                           n27105, A => n1410, ZN => n1407);
   U1566 : AOI22_X1 port map( A1 => n27101, A2 => n26701, B1 => n27097, B2 => 
                           regs_18_3_port, ZN => n1410);
   U1567 : OAI221_X1 port map( B1 => n26534, B2 => n27109, C1 => n26850, C2 => 
                           n27105, A => n1392, ZN => n1389);
   U1568 : AOI22_X1 port map( A1 => n27101, A2 => n26702, B1 => n27097, B2 => 
                           regs_18_4_port, ZN => n1392);
   U1569 : OAI221_X1 port map( B1 => n26535, B2 => n27109, C1 => n26851, C2 => 
                           n27105, A => n1374, ZN => n1371);
   U1570 : AOI22_X1 port map( A1 => n27101, A2 => n26703, B1 => n27097, B2 => 
                           regs_18_5_port, ZN => n1374);
   U1571 : OAI221_X1 port map( B1 => n26536, B2 => n27109, C1 => n26852, C2 => 
                           n27105, A => n1356, ZN => n1353);
   U1572 : AOI22_X1 port map( A1 => n27101, A2 => n26704, B1 => n27097, B2 => 
                           regs_18_6_port, ZN => n1356);
   U1573 : OAI221_X1 port map( B1 => n26537, B2 => n27109, C1 => n26853, C2 => 
                           n27105, A => n1338, ZN => n1335);
   U1574 : AOI22_X1 port map( A1 => n27101, A2 => n26705, B1 => n27097, B2 => 
                           regs_18_7_port, ZN => n1338);
   U1575 : OAI221_X1 port map( B1 => n26538, B2 => n27109, C1 => n26854, C2 => 
                           n27105, A => n1320, ZN => n1317);
   U1576 : AOI22_X1 port map( A1 => n27101, A2 => n26706, B1 => n27097, B2 => 
                           regs_18_8_port, ZN => n1320);
   U1577 : OAI221_X1 port map( B1 => n26539, B2 => n27109, C1 => n26855, C2 => 
                           n27105, A => n1292, ZN => n1283);
   U1578 : AOI22_X1 port map( A1 => n27101, A2 => n26707, B1 => n27097, B2 => 
                           regs_18_9_port, ZN => n1292);
   U1579 : OAI221_X1 port map( B1 => n26540, B2 => n27107, C1 => n26856, C2 => 
                           n27103, A => n1842, ZN => n1839);
   U1580 : AOI22_X1 port map( A1 => n27099, A2 => n26708, B1 => n27095, B2 => 
                           regs_18_10_port, ZN => n1842);
   U1581 : OAI221_X1 port map( B1 => n26541, B2 => n27107, C1 => n26857, C2 => 
                           n27103, A => n1824, ZN => n1821);
   U1582 : AOI22_X1 port map( A1 => n27099, A2 => n26709, B1 => n27095, B2 => 
                           regs_18_11_port, ZN => n1824);
   U1583 : OAI221_X1 port map( B1 => n26542, B2 => n27107, C1 => n26858, C2 => 
                           n27103, A => n1806, ZN => n1803);
   U1584 : AOI22_X1 port map( A1 => n27099, A2 => n26710, B1 => n27095, B2 => 
                           regs_18_12_port, ZN => n1806);
   U1585 : OAI221_X1 port map( B1 => n26543, B2 => n27107, C1 => n26859, C2 => 
                           n27103, A => n1788, ZN => n1785);
   U1586 : AOI22_X1 port map( A1 => n27099, A2 => n26711, B1 => n27095, B2 => 
                           regs_18_13_port, ZN => n1788);
   U1587 : OAI221_X1 port map( B1 => n26544, B2 => n27107, C1 => n26860, C2 => 
                           n27103, A => n1770, ZN => n1767);
   U1588 : AOI22_X1 port map( A1 => n27099, A2 => n26712, B1 => n27095, B2 => 
                           regs_18_14_port, ZN => n1770);
   U1589 : OAI221_X1 port map( B1 => n26545, B2 => n27107, C1 => n26861, C2 => 
                           n27103, A => n1752, ZN => n1749);
   U1590 : AOI22_X1 port map( A1 => n27099, A2 => n26713, B1 => n27095, B2 => 
                           regs_18_15_port, ZN => n1752);
   U1591 : OAI221_X1 port map( B1 => n26546, B2 => n27107, C1 => n26862, C2 => 
                           n27103, A => n1734, ZN => n1731);
   U1592 : AOI22_X1 port map( A1 => n27099, A2 => n26714, B1 => n27095, B2 => 
                           regs_18_16_port, ZN => n1734);
   U1593 : OAI221_X1 port map( B1 => n26547, B2 => n27107, C1 => n26863, C2 => 
                           n27103, A => n1716, ZN => n1713);
   U1594 : AOI22_X1 port map( A1 => n27099, A2 => n26715, B1 => n27095, B2 => 
                           regs_18_17_port, ZN => n1716);
   U1595 : OAI221_X1 port map( B1 => n26548, B2 => n27107, C1 => n26864, C2 => 
                           n27103, A => n1698, ZN => n1695);
   U1596 : AOI22_X1 port map( A1 => n27099, A2 => n26716, B1 => n27095, B2 => 
                           regs_18_18_port, ZN => n1698);
   U1597 : OAI221_X1 port map( B1 => n26549, B2 => n27107, C1 => n26865, C2 => 
                           n27103, A => n1680, ZN => n1677);
   U1598 : AOI22_X1 port map( A1 => n27099, A2 => n26717, B1 => n27095, B2 => 
                           regs_18_19_port, ZN => n1680);
   U1599 : OAI221_X1 port map( B1 => n26550, B2 => n27172, C1 => n26866, C2 => 
                           n27168, A => n1636, ZN => n1633);
   U1600 : AOI22_X1 port map( A1 => n27164, A2 => n26414, B1 => n27160, B2 => 
                           n26753, ZN => n1636);
   U1601 : OAI221_X1 port map( B1 => n26551, B2 => n27108, C1 => n26867, C2 => 
                           n27104, A => n1644, ZN => n1641);
   U1602 : AOI22_X1 port map( A1 => n27100, A2 => n26718, B1 => n27096, B2 => 
                           regs_18_20_port, ZN => n1644);
   U1603 : OAI221_X1 port map( B1 => n26552, B2 => n27172, C1 => n26868, C2 => 
                           n27168, A => n1618, ZN => n1615);
   U1604 : AOI22_X1 port map( A1 => n27164, A2 => n26415, B1 => n27160, B2 => 
                           n26754, ZN => n1618);
   U1605 : OAI221_X1 port map( B1 => n26553, B2 => n27108, C1 => n26869, C2 => 
                           n27104, A => n1626, ZN => n1623);
   U1606 : AOI22_X1 port map( A1 => n27100, A2 => n26719, B1 => n27096, B2 => 
                           regs_18_21_port, ZN => n1626);
   U1607 : OAI221_X1 port map( B1 => n26554, B2 => n27172, C1 => n26870, C2 => 
                           n27168, A => n1600, ZN => n1597);
   U1608 : AOI22_X1 port map( A1 => n27164, A2 => n26416, B1 => n27160, B2 => 
                           n26755, ZN => n1600);
   U1609 : OAI221_X1 port map( B1 => n26555, B2 => n27108, C1 => n26871, C2 => 
                           n27104, A => n1608, ZN => n1605);
   U1610 : AOI22_X1 port map( A1 => n27100, A2 => n26720, B1 => n27096, B2 => 
                           regs_18_22_port, ZN => n1608);
   U1611 : OAI221_X1 port map( B1 => n26556, B2 => n27172, C1 => n26872, C2 => 
                           n27168, A => n1582, ZN => n1579);
   U1612 : AOI22_X1 port map( A1 => n27164, A2 => n26417, B1 => n27160, B2 => 
                           n26756, ZN => n1582);
   U1613 : OAI221_X1 port map( B1 => n26557, B2 => n27108, C1 => n26873, C2 => 
                           n27104, A => n1590, ZN => n1587);
   U1614 : AOI22_X1 port map( A1 => n27100, A2 => n26721, B1 => n27096, B2 => 
                           regs_18_23_port, ZN => n1590);
   U1615 : OAI221_X1 port map( B1 => n26558, B2 => n27172, C1 => n26874, C2 => 
                           n27168, A => n1564, ZN => n1561);
   U1616 : AOI22_X1 port map( A1 => n27164, A2 => n26418, B1 => n27160, B2 => 
                           n26757, ZN => n1564);
   U1617 : OAI221_X1 port map( B1 => n26559, B2 => n27108, C1 => n26875, C2 => 
                           n27104, A => n1572, ZN => n1569);
   U1618 : AOI22_X1 port map( A1 => n27100, A2 => n26722, B1 => n27096, B2 => 
                           regs_18_24_port, ZN => n1572);
   U1619 : OAI221_X1 port map( B1 => n26560, B2 => n27172, C1 => n26876, C2 => 
                           n27168, A => n1546, ZN => n1543);
   U1620 : AOI22_X1 port map( A1 => n27164, A2 => n26419, B1 => n27160, B2 => 
                           n26758, ZN => n1546);
   U1621 : OAI221_X1 port map( B1 => n26561, B2 => n27108, C1 => n26877, C2 => 
                           n27104, A => n1554, ZN => n1551);
   U1622 : AOI22_X1 port map( A1 => n27100, A2 => n26723, B1 => n27096, B2 => 
                           regs_18_25_port, ZN => n1554);
   U1623 : OAI221_X1 port map( B1 => n26562, B2 => n27172, C1 => n26878, C2 => 
                           n27168, A => n1528, ZN => n1525);
   U1624 : AOI22_X1 port map( A1 => n27164, A2 => n26420, B1 => n27160, B2 => 
                           n26759, ZN => n1528);
   U1625 : OAI221_X1 port map( B1 => n26563, B2 => n27108, C1 => n26879, C2 => 
                           n27104, A => n1536, ZN => n1533);
   U1626 : AOI22_X1 port map( A1 => n27100, A2 => n26724, B1 => n27096, B2 => 
                           regs_18_26_port, ZN => n1536);
   U1627 : OAI221_X1 port map( B1 => n26564, B2 => n27172, C1 => n26880, C2 => 
                           n27168, A => n1510, ZN => n1507);
   U1628 : AOI22_X1 port map( A1 => n27164, A2 => n26421, B1 => n27160, B2 => 
                           n26760, ZN => n1510);
   U1629 : OAI221_X1 port map( B1 => n26565, B2 => n27108, C1 => n26881, C2 => 
                           n27104, A => n1518, ZN => n1515);
   U1630 : AOI22_X1 port map( A1 => n27100, A2 => n26725, B1 => n27096, B2 => 
                           regs_18_27_port, ZN => n1518);
   U1631 : OAI221_X1 port map( B1 => n26566, B2 => n27172, C1 => n26882, C2 => 
                           n27168, A => n1492, ZN => n1489);
   U1632 : AOI22_X1 port map( A1 => n27164, A2 => n26422, B1 => n27160, B2 => 
                           n26761, ZN => n1492);
   U1633 : OAI221_X1 port map( B1 => n26567, B2 => n27108, C1 => n26883, C2 => 
                           n27104, A => n1500, ZN => n1497);
   U1634 : AOI22_X1 port map( A1 => n27100, A2 => n26726, B1 => n27096, B2 => 
                           regs_18_28_port, ZN => n1500);
   U1635 : OAI221_X1 port map( B1 => n26568, B2 => n27172, C1 => n26884, C2 => 
                           n27168, A => n1474, ZN => n1471);
   U1636 : AOI22_X1 port map( A1 => n27164, A2 => n26423, B1 => n27160, B2 => 
                           n26762, ZN => n1474);
   U1637 : OAI221_X1 port map( B1 => n26569, B2 => n27108, C1 => n26885, C2 => 
                           n27104, A => n1482, ZN => n1479);
   U1638 : AOI22_X1 port map( A1 => n27100, A2 => n26727, B1 => n27096, B2 => 
                           regs_18_29_port, ZN => n1482);
   U1639 : OAI221_X1 port map( B1 => n26570, B2 => n27173, C1 => n26886, C2 => 
                           n27169, A => n1438, ZN => n1435);
   U1640 : AOI22_X1 port map( A1 => n27165, A2 => n26424, B1 => n27161, B2 => 
                           n26763, ZN => n1438);
   U1641 : OAI221_X1 port map( B1 => n26571, B2 => n27109, C1 => n26887, C2 => 
                           n27105, A => n1446, ZN => n1443);
   U1642 : AOI22_X1 port map( A1 => n27101, A2 => n26728, B1 => n27097, B2 => 
                           regs_18_30_port, ZN => n1446);
   U1643 : OAI221_X1 port map( B1 => n26572, B2 => n27173, C1 => n26888, C2 => 
                           n27169, A => n1420, ZN => n1417);
   U1644 : AOI22_X1 port map( A1 => n27165, A2 => n26425, B1 => n27161, B2 => 
                           n26764, ZN => n1420);
   U1645 : OAI221_X1 port map( B1 => n26573, B2 => n27109, C1 => n26889, C2 => 
                           n27105, A => n1428, ZN => n1425);
   U1646 : AOI22_X1 port map( A1 => n27101, A2 => n26729, B1 => n27097, B2 => 
                           regs_18_31_port, ZN => n1428);
   U1647 : OAI221_X1 port map( B1 => n25511, B2 => n27091, C1 => n26596, C2 => 
                           n27087, A => n1825, ZN => n1820);
   U1648 : AOI22_X1 port map( A1 => n27083, A2 => n25445, B1 => n27079, B2 => 
                           n26589, ZN => n1825);
   U1649 : OAI221_X1 port map( B1 => n25512, B2 => n27091, C1 => n26597, C2 => 
                           n27087, A => n1807, ZN => n1802);
   U1650 : AOI22_X1 port map( A1 => n27083, A2 => n25446, B1 => n27079, B2 => 
                           n26590, ZN => n1807);
   U1651 : OAI221_X1 port map( B1 => n25513, B2 => n27091, C1 => n26598, C2 => 
                           n27087, A => n1789, ZN => n1784);
   U1652 : AOI22_X1 port map( A1 => n27083, A2 => n25447, B1 => n27079, B2 => 
                           n26591, ZN => n1789);
   U1653 : OAI221_X1 port map( B1 => n25514, B2 => n27091, C1 => n26599, C2 => 
                           n27087, A => n1771, ZN => n1766);
   U1654 : AOI22_X1 port map( A1 => n27083, A2 => n25448, B1 => n27079, B2 => 
                           n26592, ZN => n1771);
   U1655 : OAI221_X1 port map( B1 => n25532, B2 => n26964, C1 => n25291, C2 => 
                           n26967, A => n1253, ZN => n1246);
   U1656 : AOI22_X1 port map( A1 => n25211, A2 => n27710, B1 => n25466, B2 => 
                           n27711, ZN => n1253);
   U1657 : OAI221_X1 port map( B1 => n25533, B2 => n26966, C1 => n25292, C2 => 
                           n26969, A => n1043_port, ZN => n1038_port);
   U1658 : AOI22_X1 port map( A1 => n25212, A2 => n27710, B1 => n25467, B2 => 
                           n27711, ZN => n1043_port);
   U1659 : OAI221_X1 port map( B1 => n25534, B2 => n26966, C1 => n25293, C2 => 
                           n26969, A => n845_port, ZN => n840_port);
   U1660 : AOI22_X1 port map( A1 => n25213, A2 => n27710, B1 => n25468, B2 => 
                           n27711, ZN => n845_port);
   U1661 : OAI221_X1 port map( B1 => n25535, B2 => n26964, C1 => n25294, C2 => 
                           n26967, A => n785_port, ZN => n780_port);
   U1662 : AOI22_X1 port map( A1 => n25214, A2 => n27710, B1 => n25469, B2 => 
                           n27711, ZN => n785_port);
   U1663 : OAI221_X1 port map( B1 => n25536, B2 => n26964, C1 => n25295, C2 => 
                           n26967, A => n767_port, ZN => n762_port);
   U1664 : AOI22_X1 port map( A1 => n25215, A2 => n27710, B1 => n25470, B2 => 
                           n27711, ZN => n767_port);
   U1665 : OAI221_X1 port map( B1 => n25537, B2 => n26965, C1 => n25296, C2 => 
                           n26968, A => n749_port, ZN => n744_port);
   U1666 : AOI22_X1 port map( A1 => n25216, A2 => n27710, B1 => n25471, B2 => 
                           n27711, ZN => n749_port);
   U1667 : OAI221_X1 port map( B1 => n25538, B2 => n26966, C1 => n25297, C2 => 
                           n26969, A => n731_port, ZN => n726_port);
   U1668 : AOI22_X1 port map( A1 => n25217, A2 => n27710, B1 => n25472, B2 => 
                           n27711, ZN => n731_port);
   U1669 : OAI221_X1 port map( B1 => n25539, B2 => n26965, C1 => n25298, C2 => 
                           n26968, A => n713_port, ZN => n708_port);
   U1670 : AOI22_X1 port map( A1 => n25218, A2 => n27710, B1 => n25473, B2 => 
                           n27711, ZN => n713_port);
   U1671 : OAI221_X1 port map( B1 => n25540, B2 => n26964, C1 => n25299, C2 => 
                           n26967, A => n695_port, ZN => n690_port);
   U1672 : AOI22_X1 port map( A1 => n25219, A2 => n27710, B1 => n25474, B2 => 
                           n27711, ZN => n695_port);
   U1673 : OAI221_X1 port map( B1 => n25541, B2 => n26965, C1 => n25300, C2 => 
                           n26968, A => n675_port, ZN => n660_port);
   U1674 : AOI22_X1 port map( A1 => n25220, A2 => n27710, B1 => n25475, B2 => 
                           n27711, ZN => n675_port);
   U1675 : OAI221_X1 port map( B1 => n25542, B2 => n26965, C1 => n25301, C2 => 
                           n26968, A => n1223, ZN => n1218);
   U1676 : AOI22_X1 port map( A1 => n25221, A2 => n27710, B1 => n25476, B2 => 
                           n27711, ZN => n1223);
   U1677 : OAI221_X1 port map( B1 => n25543, B2 => n26966, C1 => n25302, C2 => 
                           n26969, A => n1205, ZN => n1200);
   U1678 : AOI22_X1 port map( A1 => n25222, A2 => n27710, B1 => n25477, B2 => 
                           n27711, ZN => n1205);
   U1679 : OAI221_X1 port map( B1 => n25544, B2 => n26966, C1 => n25303, C2 => 
                           n26969, A => n1187, ZN => n1182);
   U1680 : AOI22_X1 port map( A1 => n25223, A2 => n27710, B1 => n25478, B2 => 
                           n27711, ZN => n1187);
   U1681 : OAI221_X1 port map( B1 => n25545, B2 => n26964, C1 => n25304, C2 => 
                           n26967, A => n1169, ZN => n1164);
   U1682 : AOI22_X1 port map( A1 => n25224, A2 => n27710, B1 => n25479, B2 => 
                           n27711, ZN => n1169);
   U1683 : OAI221_X1 port map( B1 => n25546, B2 => n26964, C1 => n25305, C2 => 
                           n26967, A => n1151, ZN => n1146);
   U1684 : AOI22_X1 port map( A1 => n25225, A2 => n27710, B1 => n25480, B2 => 
                           n27711, ZN => n1151);
   U1685 : OAI221_X1 port map( B1 => n25547, B2 => n26965, C1 => n25306, C2 => 
                           n26968, A => n1133, ZN => n1128);
   U1686 : AOI22_X1 port map( A1 => n25226, A2 => n27710, B1 => n25481, B2 => 
                           n27711, ZN => n1133);
   U1687 : OAI221_X1 port map( B1 => n25548, B2 => n26966, C1 => n25307, C2 => 
                           n26969, A => n1115, ZN => n1110);
   U1688 : AOI22_X1 port map( A1 => n25227, A2 => n27710, B1 => n25482, B2 => 
                           n27711, ZN => n1115);
   U1689 : OAI221_X1 port map( B1 => n25549, B2 => n26965, C1 => n25308, C2 => 
                           n26968, A => n1097, ZN => n1092);
   U1690 : AOI22_X1 port map( A1 => n25228, A2 => n27710, B1 => n25483, B2 => 
                           n27711, ZN => n1097);
   U1691 : OAI221_X1 port map( B1 => n25550, B2 => n26964, C1 => n25309, C2 => 
                           n26967, A => n1079, ZN => n1074);
   U1692 : AOI22_X1 port map( A1 => n25229, A2 => n27710, B1 => n25484, B2 => 
                           n27711, ZN => n1079);
   U1693 : OAI221_X1 port map( B1 => n25551, B2 => n26965, C1 => n25310, C2 => 
                           n26968, A => n1061, ZN => n1056);
   U1694 : AOI22_X1 port map( A1 => n25230, A2 => n27710, B1 => n25485, B2 => 
                           n27711, ZN => n1061);
   U1695 : OAI221_X1 port map( B1 => n25500, B2 => n27091, C1 => n25259, C2 => 
                           n27087, A => n1873, ZN => n1866);
   U1696 : AOI22_X1 port map( A1 => n27083, A2 => n25434, B1 => n27079, B2 => 
                           n25179, ZN => n1873);
   U1697 : OAI221_X1 port map( B1 => n25501, B2 => n27092, C1 => n25260, C2 => 
                           n27088, A => n1663, ZN => n1658);
   U1698 : AOI22_X1 port map( A1 => n27084, A2 => n25435, B1 => n27080, B2 => 
                           n25180, ZN => n1663);
   U1699 : OAI221_X1 port map( B1 => n25502, B2 => n27093, C1 => n25261, C2 => 
                           n27089, A => n1465, ZN => n1460);
   U1700 : AOI22_X1 port map( A1 => n27085, A2 => n25436, B1 => n27081, B2 => 
                           n25181, ZN => n1465);
   U1701 : OAI221_X1 port map( B1 => n25503, B2 => n27093, C1 => n25262, C2 => 
                           n27089, A => n1411, ZN => n1406);
   U1702 : AOI22_X1 port map( A1 => n27085, A2 => n25437, B1 => n27081, B2 => 
                           n25182, ZN => n1411);
   U1703 : OAI221_X1 port map( B1 => n25504, B2 => n27093, C1 => n25263, C2 => 
                           n27089, A => n1393, ZN => n1388);
   U1704 : AOI22_X1 port map( A1 => n27085, A2 => n25438, B1 => n27081, B2 => 
                           n25183, ZN => n1393);
   U1705 : OAI221_X1 port map( B1 => n25505, B2 => n27093, C1 => n25264, C2 => 
                           n27089, A => n1375, ZN => n1370);
   U1706 : AOI22_X1 port map( A1 => n27085, A2 => n25439, B1 => n27081, B2 => 
                           n25184, ZN => n1375);
   U1707 : OAI221_X1 port map( B1 => n25506, B2 => n27093, C1 => n25265, C2 => 
                           n27089, A => n1357, ZN => n1352);
   U1708 : AOI22_X1 port map( A1 => n27085, A2 => n25440, B1 => n27081, B2 => 
                           n25185, ZN => n1357);
   U1709 : OAI221_X1 port map( B1 => n25507, B2 => n27093, C1 => n25266, C2 => 
                           n27089, A => n1339, ZN => n1334);
   U1710 : AOI22_X1 port map( A1 => n27085, A2 => n25441, B1 => n27081, B2 => 
                           n25186, ZN => n1339);
   U1711 : OAI221_X1 port map( B1 => n25508, B2 => n27093, C1 => n25267, C2 => 
                           n27089, A => n1321, ZN => n1316);
   U1712 : AOI22_X1 port map( A1 => n27085, A2 => n25442, B1 => n27081, B2 => 
                           n26593, ZN => n1321);
   U1713 : OAI221_X1 port map( B1 => n25509, B2 => n27093, C1 => n25268, C2 => 
                           n27089, A => n1297, ZN => n1282);
   U1714 : AOI22_X1 port map( A1 => n27085, A2 => n25443, B1 => n27081, B2 => 
                           n26594, ZN => n1297);
   U1715 : OAI221_X1 port map( B1 => n25510, B2 => n27091, C1 => n25269, C2 => 
                           n27087, A => n1843, ZN => n1838);
   U1716 : AOI22_X1 port map( A1 => n27083, A2 => n25444, B1 => n27079, B2 => 
                           n26595, ZN => n1843);
   U1717 : OAI221_X1 port map( B1 => n25515, B2 => n27091, C1 => n26890, C2 => 
                           n27087, A => n1753, ZN => n1748);
   U1718 : AOI22_X1 port map( A1 => n27083, A2 => n26426, B1 => n27079, B2 => 
                           n26765, ZN => n1753);
   U1719 : OAI221_X1 port map( B1 => n25516, B2 => n27091, C1 => n26891, C2 => 
                           n27087, A => n1735, ZN => n1730);
   U1720 : AOI22_X1 port map( A1 => n27083, A2 => n26427, B1 => n27079, B2 => 
                           n26766, ZN => n1735);
   U1721 : OAI221_X1 port map( B1 => n26327, B2 => n27155, C1 => n26600, C2 => 
                           n27151, A => n1859, ZN => n1848);
   U1722 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_0_port, B1 => n27143, 
                           B2 => regs_13_0_port, ZN => n1859);
   U1723 : OAI221_X1 port map( B1 => n26328, B2 => n27156, C1 => n26601, C2 => 
                           n27152, A => n1655, ZN => n1650);
   U1724 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_1_port, B1 => n27144, 
                           B2 => regs_13_1_port, ZN => n1655);
   U1725 : OAI221_X1 port map( B1 => n26329, B2 => n27157, C1 => n26602, C2 => 
                           n27153, A => n1457, ZN => n1452);
   U1726 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_2_port, B1 => n27145, 
                           B2 => regs_13_2_port, ZN => n1457);
   U1727 : OAI221_X1 port map( B1 => n26330, B2 => n27157, C1 => n26603, C2 => 
                           n27153, A => n1403, ZN => n1398);
   U1728 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_3_port, B1 => n27145, 
                           B2 => regs_13_3_port, ZN => n1403);
   U1729 : OAI221_X1 port map( B1 => n26331, B2 => n27157, C1 => n26604, C2 => 
                           n27153, A => n1385, ZN => n1380);
   U1730 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_4_port, B1 => n27145, 
                           B2 => regs_13_4_port, ZN => n1385);
   U1731 : OAI221_X1 port map( B1 => n26332, B2 => n27157, C1 => n26605, C2 => 
                           n27153, A => n1367, ZN => n1362);
   U1732 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_5_port, B1 => n27145, 
                           B2 => regs_13_5_port, ZN => n1367);
   U1733 : OAI221_X1 port map( B1 => n26333, B2 => n27157, C1 => n26606, C2 => 
                           n27153, A => n1349, ZN => n1344);
   U1734 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_6_port, B1 => n27145, 
                           B2 => regs_13_6_port, ZN => n1349);
   U1735 : OAI221_X1 port map( B1 => n26334, B2 => n27157, C1 => n26607, C2 => 
                           n27153, A => n1331, ZN => n1326);
   U1736 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_7_port, B1 => n27145, 
                           B2 => regs_13_7_port, ZN => n1331);
   U1737 : OAI221_X1 port map( B1 => n26335, B2 => n27157, C1 => n26608, C2 => 
                           n27153, A => n1313, ZN => n1308);
   U1738 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_8_port, B1 => n27145, 
                           B2 => regs_13_8_port, ZN => n1313);
   U1739 : OAI221_X1 port map( B1 => n26336, B2 => n27157, C1 => n26609, C2 => 
                           n27153, A => n1273, ZN => n1258);
   U1740 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_9_port, B1 => n27145, 
                           B2 => regs_13_9_port, ZN => n1273);
   U1741 : OAI221_X1 port map( B1 => n26337, B2 => n27155, C1 => n26610, C2 => 
                           n27151, A => n1835, ZN => n1830);
   U1742 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_10_port, B1 => n27143,
                           B2 => regs_13_10_port, ZN => n1835);
   U1743 : OAI221_X1 port map( B1 => n26338, B2 => n27155, C1 => n26611, C2 => 
                           n27151, A => n1817, ZN => n1812);
   U1744 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_11_port, B1 => n27143,
                           B2 => regs_13_11_port, ZN => n1817);
   U1745 : OAI221_X1 port map( B1 => n26339, B2 => n27155, C1 => n26612, C2 => 
                           n27151, A => n1799, ZN => n1794);
   U1746 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_12_port, B1 => n27143,
                           B2 => regs_13_12_port, ZN => n1799);
   U1747 : OAI221_X1 port map( B1 => n26340, B2 => n27155, C1 => n26613, C2 => 
                           n27151, A => n1781, ZN => n1776);
   U1748 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_13_port, B1 => n27143,
                           B2 => regs_13_13_port, ZN => n1781);
   U1749 : OAI221_X1 port map( B1 => n26341, B2 => n27155, C1 => n26614, C2 => 
                           n27151, A => n1763, ZN => n1758);
   U1750 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_14_port, B1 => n27143,
                           B2 => regs_13_14_port, ZN => n1763);
   U1751 : OAI221_X1 port map( B1 => n26342, B2 => n27155, C1 => n26615, C2 => 
                           n27151, A => n1745, ZN => n1740);
   U1752 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_15_port, B1 => n27143,
                           B2 => regs_13_15_port, ZN => n1745);
   U1753 : OAI221_X1 port map( B1 => n26343, B2 => n27155, C1 => n26616, C2 => 
                           n27151, A => n1727, ZN => n1722);
   U1754 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_16_port, B1 => n27143,
                           B2 => regs_13_16_port, ZN => n1727);
   U1755 : OAI221_X1 port map( B1 => n26344, B2 => n27155, C1 => n26617, C2 => 
                           n27151, A => n1709, ZN => n1704);
   U1756 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_17_port, B1 => n27143,
                           B2 => regs_13_17_port, ZN => n1709);
   U1757 : OAI221_X1 port map( B1 => n26574, B2 => n27091, C1 => n26892, C2 => 
                           n27087, A => n1717, ZN => n1712);
   U1758 : AOI22_X1 port map( A1 => n27083, A2 => n26428, B1 => n27079, B2 => 
                           n26767, ZN => n1717);
   U1759 : OAI221_X1 port map( B1 => n26345, B2 => n27155, C1 => n26618, C2 => 
                           n27151, A => n1691, ZN => n1686);
   U1760 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_18_port, B1 => n27143,
                           B2 => regs_13_18_port, ZN => n1691);
   U1761 : OAI221_X1 port map( B1 => n26575, B2 => n27091, C1 => n26893, C2 => 
                           n27087, A => n1699, ZN => n1694);
   U1762 : AOI22_X1 port map( A1 => n27083, A2 => n26429, B1 => n27079, B2 => 
                           n26768, ZN => n1699);
   U1763 : OAI221_X1 port map( B1 => n26346, B2 => n27155, C1 => n26619, C2 => 
                           n27151, A => n1673, ZN => n1668);
   U1764 : AOI22_X1 port map( A1 => n27147, A2 => regs_5_19_port, B1 => n27143,
                           B2 => regs_13_19_port, ZN => n1673);
   U1765 : OAI221_X1 port map( B1 => n26576, B2 => n27091, C1 => n26894, C2 => 
                           n27087, A => n1681, ZN => n1676);
   U1766 : AOI22_X1 port map( A1 => n27083, A2 => n26430, B1 => n27079, B2 => 
                           n26769, ZN => n1681);
   U1767 : OAI221_X1 port map( B1 => n26347, B2 => n27156, C1 => n26620, C2 => 
                           n27152, A => n1637, ZN => n1632);
   U1768 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_20_port, B1 => n27144,
                           B2 => regs_13_20_port, ZN => n1637);
   U1769 : OAI221_X1 port map( B1 => n26577, B2 => n27092, C1 => n26895, C2 => 
                           n27088, A => n1645, ZN => n1640);
   U1770 : AOI22_X1 port map( A1 => n27084, A2 => n26431, B1 => n27080, B2 => 
                           n26770, ZN => n1645);
   U1771 : OAI221_X1 port map( B1 => n26348, B2 => n27156, C1 => n26621, C2 => 
                           n27152, A => n1619, ZN => n1614);
   U1772 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_21_port, B1 => n27144,
                           B2 => regs_13_21_port, ZN => n1619);
   U1773 : OAI221_X1 port map( B1 => n26578, B2 => n27092, C1 => n26896, C2 => 
                           n27088, A => n1627, ZN => n1622);
   U1774 : AOI22_X1 port map( A1 => n27084, A2 => n26432, B1 => n27080, B2 => 
                           n26771, ZN => n1627);
   U1775 : OAI221_X1 port map( B1 => n26349, B2 => n27156, C1 => n26622, C2 => 
                           n27152, A => n1601, ZN => n1596);
   U1776 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_22_port, B1 => n27144,
                           B2 => regs_13_22_port, ZN => n1601);
   U1777 : OAI221_X1 port map( B1 => n26579, B2 => n27092, C1 => n26897, C2 => 
                           n27088, A => n1609, ZN => n1604);
   U1778 : AOI22_X1 port map( A1 => n27084, A2 => n26433, B1 => n27080, B2 => 
                           n26772, ZN => n1609);
   U1779 : OAI221_X1 port map( B1 => n26350, B2 => n27156, C1 => n26623, C2 => 
                           n27152, A => n1583, ZN => n1578);
   U1780 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_23_port, B1 => n27144,
                           B2 => regs_13_23_port, ZN => n1583);
   U1781 : OAI221_X1 port map( B1 => n26580, B2 => n27092, C1 => n26898, C2 => 
                           n27088, A => n1591, ZN => n1586);
   U1782 : AOI22_X1 port map( A1 => n27084, A2 => n26434, B1 => n27080, B2 => 
                           n26773, ZN => n1591);
   U1783 : OAI221_X1 port map( B1 => n26351, B2 => n27156, C1 => n26624, C2 => 
                           n27152, A => n1565, ZN => n1560);
   U1784 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_24_port, B1 => n27144,
                           B2 => regs_13_24_port, ZN => n1565);
   U1785 : OAI221_X1 port map( B1 => n26581, B2 => n27092, C1 => n26899, C2 => 
                           n27088, A => n1573, ZN => n1568);
   U1786 : AOI22_X1 port map( A1 => n27084, A2 => n26435, B1 => n27080, B2 => 
                           n26774, ZN => n1573);
   U1787 : OAI221_X1 port map( B1 => n26352, B2 => n27156, C1 => n26625, C2 => 
                           n27152, A => n1547, ZN => n1542);
   U1788 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_25_port, B1 => n27144,
                           B2 => regs_13_25_port, ZN => n1547);
   U1789 : OAI221_X1 port map( B1 => n26582, B2 => n27092, C1 => n26900, C2 => 
                           n27088, A => n1555, ZN => n1550);
   U1790 : AOI22_X1 port map( A1 => n27084, A2 => n26436, B1 => n27080, B2 => 
                           n26775, ZN => n1555);
   U1791 : OAI221_X1 port map( B1 => n26353, B2 => n27156, C1 => n26626, C2 => 
                           n27152, A => n1529, ZN => n1524);
   U1792 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_26_port, B1 => n27144,
                           B2 => regs_13_26_port, ZN => n1529);
   U1793 : OAI221_X1 port map( B1 => n26583, B2 => n27092, C1 => n26901, C2 => 
                           n27088, A => n1537, ZN => n1532);
   U1794 : AOI22_X1 port map( A1 => n27084, A2 => n26437, B1 => n27080, B2 => 
                           n26776, ZN => n1537);
   U1795 : OAI221_X1 port map( B1 => n26354, B2 => n27156, C1 => n26627, C2 => 
                           n27152, A => n1511, ZN => n1506);
   U1796 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_27_port, B1 => n27144,
                           B2 => regs_13_27_port, ZN => n1511);
   U1797 : OAI221_X1 port map( B1 => n26584, B2 => n27092, C1 => n26902, C2 => 
                           n27088, A => n1519, ZN => n1514);
   U1798 : AOI22_X1 port map( A1 => n27084, A2 => n26438, B1 => n27080, B2 => 
                           n26777, ZN => n1519);
   U1799 : OAI221_X1 port map( B1 => n26355, B2 => n27156, C1 => n26628, C2 => 
                           n27152, A => n1493, ZN => n1488);
   U1800 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_28_port, B1 => n27144,
                           B2 => regs_13_28_port, ZN => n1493);
   U1801 : OAI221_X1 port map( B1 => n26585, B2 => n27092, C1 => n26903, C2 => 
                           n27088, A => n1501, ZN => n1496);
   U1802 : AOI22_X1 port map( A1 => n27084, A2 => n26439, B1 => n27080, B2 => 
                           n26778, ZN => n1501);
   U1803 : OAI221_X1 port map( B1 => n26356, B2 => n27156, C1 => n26629, C2 => 
                           n27152, A => n1475, ZN => n1470);
   U1804 : AOI22_X1 port map( A1 => n27148, A2 => regs_5_29_port, B1 => n27144,
                           B2 => regs_13_29_port, ZN => n1475);
   U1805 : OAI221_X1 port map( B1 => n26586, B2 => n27092, C1 => n26904, C2 => 
                           n27088, A => n1483, ZN => n1478);
   U1806 : AOI22_X1 port map( A1 => n27084, A2 => n26440, B1 => n27080, B2 => 
                           n26779, ZN => n1483);
   U1807 : OAI221_X1 port map( B1 => n26357, B2 => n27157, C1 => n26630, C2 => 
                           n27153, A => n1439, ZN => n1434);
   U1808 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_30_port, B1 => n27145,
                           B2 => regs_13_30_port, ZN => n1439);
   U1809 : OAI221_X1 port map( B1 => n26587, B2 => n27093, C1 => n26905, C2 => 
                           n27089, A => n1447, ZN => n1442);
   U1810 : AOI22_X1 port map( A1 => n27085, A2 => n26441, B1 => n27081, B2 => 
                           n26780, ZN => n1447);
   U1811 : OAI221_X1 port map( B1 => n26358, B2 => n27157, C1 => n26631, C2 => 
                           n27153, A => n1421, ZN => n1416);
   U1812 : AOI22_X1 port map( A1 => n27149, A2 => regs_5_31_port, B1 => n27145,
                           B2 => regs_13_31_port, ZN => n1421);
   U1813 : OAI221_X1 port map( B1 => n26588, B2 => n27093, C1 => n26906, C2 => 
                           n27089, A => n1429, ZN => n1424);
   U1814 : AOI22_X1 port map( A1 => n27085, A2 => n26442, B1 => n27081, B2 => 
                           n26781, ZN => n1429);
   U1815 : AND2_X1 port map( A1 => add_rd2(4), A2 => n27714, ZN => n1240);
   U1816 : OAI221_X1 port map( B1 => n1889, B2 => n27241, C1 => n1890, C2 => 
                           n27237, A => n1244, ZN => n1227);
   U1817 : AOI22_X1 port map( A1 => n1887, A2 => n27233, B1 => n1888, B2 => 
                           n27229, ZN => n1244);
   U1818 : OAI221_X1 port map( B1 => n1893, B2 => n27242, C1 => n1894, C2 => 
                           n27238, A => n1036_port, ZN => n1029_port);
   U1819 : AOI22_X1 port map( A1 => n1891, A2 => n27233, B1 => n1892, B2 => 
                           n27229, ZN => n1036_port);
   U1820 : OAI221_X1 port map( B1 => n1897, B2 => n27243, C1 => n1898, C2 => 
                           n27239, A => n838_port, ZN => n831_port);
   U1821 : AOI22_X1 port map( A1 => n1895, A2 => n27234, B1 => n1896, B2 => 
                           n27230, ZN => n838_port);
   U1822 : OAI221_X1 port map( B1 => n1901, B2 => n27243, C1 => n1902, C2 => 
                           n27239, A => n778_port, ZN => n771_port);
   U1823 : AOI22_X1 port map( A1 => n1899, A2 => n27235, B1 => n1900, B2 => 
                           n27231, ZN => n778_port);
   U1824 : OAI221_X1 port map( B1 => n1905, B2 => n27243, C1 => n1906, C2 => 
                           n27239, A => n760_port, ZN => n753_port);
   U1825 : AOI22_X1 port map( A1 => n1903, A2 => n27235, B1 => n1904, B2 => 
                           n27231, ZN => n760_port);
   U1826 : OAI221_X1 port map( B1 => n1909, B2 => n27243, C1 => n1910, C2 => 
                           n27239, A => n742_port, ZN => n735_port);
   U1827 : AOI22_X1 port map( A1 => n1907, A2 => n27235, B1 => n1908, B2 => 
                           n27231, ZN => n742_port);
   U1828 : OAI221_X1 port map( B1 => n1913, B2 => n27243, C1 => n1914, C2 => 
                           n27239, A => n724_port, ZN => n717_port);
   U1829 : AOI22_X1 port map( A1 => n1911, A2 => n27235, B1 => n1912, B2 => 
                           n27231, ZN => n724_port);
   U1830 : OAI221_X1 port map( B1 => n1917, B2 => n27243, C1 => n1918, C2 => 
                           n27239, A => n706_port, ZN => n699_port);
   U1831 : AOI22_X1 port map( A1 => n1915, A2 => n27235, B1 => n1916, B2 => 
                           n27231, ZN => n706_port);
   U1832 : OAI221_X1 port map( B1 => n1921, B2 => n27243, C1 => n1922, C2 => 
                           n27239, A => n688_port, ZN => n681_port);
   U1833 : AOI22_X1 port map( A1 => n1919, A2 => n27235, B1 => n1920, B2 => 
                           n27231, ZN => n688_port);
   U1834 : OAI221_X1 port map( B1 => n1925, B2 => n27243, C1 => n1926, C2 => 
                           n27239, A => n656_port, ZN => n637_port);
   U1835 : AOI22_X1 port map( A1 => n1923, A2 => n27235, B1 => n1924, B2 => 
                           n27231, ZN => n656_port);
   U1836 : OAI221_X1 port map( B1 => n1929, B2 => n27241, C1 => n1930, C2 => 
                           n27237, A => n1216, ZN => n1209);
   U1837 : AOI22_X1 port map( A1 => n1927, A2 => n27233, B1 => n1928, B2 => 
                           n27229, ZN => n1216);
   U1838 : OAI221_X1 port map( B1 => n1933, B2 => n27241, C1 => n1934, C2 => 
                           n27237, A => n1198, ZN => n1191);
   U1839 : AOI22_X1 port map( A1 => n1931, A2 => n27233, B1 => n1932, B2 => 
                           n27229, ZN => n1198);
   U1840 : OAI221_X1 port map( B1 => n1937, B2 => n27241, C1 => n1938, C2 => 
                           n27237, A => n1180, ZN => n1173);
   U1841 : AOI22_X1 port map( A1 => n1935, A2 => n27233, B1 => n1936, B2 => 
                           n27229, ZN => n1180);
   U1842 : OAI221_X1 port map( B1 => n1941, B2 => n27241, C1 => n1942, C2 => 
                           n27237, A => n1162, ZN => n1155);
   U1843 : AOI22_X1 port map( A1 => n1939, A2 => n27233, B1 => n1940, B2 => 
                           n27229, ZN => n1162);
   U1844 : OAI221_X1 port map( B1 => n1945, B2 => n27241, C1 => n1946, C2 => 
                           n27237, A => n1144, ZN => n1137);
   U1845 : AOI22_X1 port map( A1 => n1943, A2 => n27233, B1 => n1944, B2 => 
                           n27229, ZN => n1144);
   U1846 : OAI221_X1 port map( B1 => n1949, B2 => n27241, C1 => n1950, C2 => 
                           n27237, A => n1126, ZN => n1119);
   U1847 : AOI22_X1 port map( A1 => n1947, A2 => n27233, B1 => n1948, B2 => 
                           n27229, ZN => n1126);
   U1848 : OAI221_X1 port map( B1 => n1953, B2 => n27241, C1 => n1954, C2 => 
                           n27237, A => n1108, ZN => n1101);
   U1849 : AOI22_X1 port map( A1 => n1951, A2 => n27233, B1 => n1952, B2 => 
                           n27229, ZN => n1108);
   U1850 : OAI221_X1 port map( B1 => n1957, B2 => n27241, C1 => n1958, C2 => 
                           n27237, A => n1090, ZN => n1083);
   U1851 : AOI22_X1 port map( A1 => n1955, A2 => n27233, B1 => n1956, B2 => 
                           n27229, ZN => n1090);
   U1852 : OAI221_X1 port map( B1 => n1961, B2 => n27241, C1 => n1962, C2 => 
                           n27237, A => n1072, ZN => n1065);
   U1853 : AOI22_X1 port map( A1 => n1959, A2 => n27233, B1 => n1960, B2 => 
                           n27229, ZN => n1072);
   U1854 : OAI221_X1 port map( B1 => n1965, B2 => n27241, C1 => n1966, C2 => 
                           n27237, A => n1054, ZN => n1047);
   U1855 : AOI22_X1 port map( A1 => n1963, A2 => n27233, B1 => n1964, B2 => 
                           n27229, ZN => n1054);
   U1856 : OAI221_X1 port map( B1 => n1969, B2 => n27242, C1 => n1970, C2 => 
                           n27238, A => n1018_port, ZN => n1011_port);
   U1857 : AOI22_X1 port map( A1 => n1967, A2 => n27234, B1 => n1968, B2 => 
                           n27230, ZN => n1018_port);
   U1858 : OAI221_X1 port map( B1 => n1973, B2 => n27242, C1 => n1974, C2 => 
                           n27238, A => n1000_port, ZN => n993_port);
   U1859 : AOI22_X1 port map( A1 => n1971, A2 => n27234, B1 => n1972, B2 => 
                           n27230, ZN => n1000_port);
   U1860 : OAI221_X1 port map( B1 => n1977, B2 => n27242, C1 => n1978, C2 => 
                           n27238, A => n982_port, ZN => n975_port);
   U1861 : AOI22_X1 port map( A1 => n1975, A2 => n27234, B1 => n1976, B2 => 
                           n27230, ZN => n982_port);
   U1862 : OAI221_X1 port map( B1 => n1981, B2 => n27242, C1 => n1982, C2 => 
                           n27238, A => n964_port, ZN => n957_port);
   U1863 : AOI22_X1 port map( A1 => n1979, A2 => n27234, B1 => n1980, B2 => 
                           n27230, ZN => n964_port);
   U1864 : OAI221_X1 port map( B1 => n1985, B2 => n27242, C1 => n1986, C2 => 
                           n27238, A => n946_port, ZN => n939_port);
   U1865 : AOI22_X1 port map( A1 => n1983, A2 => n27234, B1 => n1984, B2 => 
                           n27230, ZN => n946_port);
   U1866 : OAI221_X1 port map( B1 => n1989, B2 => n27242, C1 => n1990, C2 => 
                           n27238, A => n928_port, ZN => n921_port);
   U1867 : AOI22_X1 port map( A1 => n1987, A2 => n27234, B1 => n1988, B2 => 
                           n27230, ZN => n928_port);
   U1868 : OAI221_X1 port map( B1 => n1993, B2 => n27242, C1 => n1994, C2 => 
                           n27238, A => n910_port, ZN => n903_port);
   U1869 : AOI22_X1 port map( A1 => n1991, A2 => n27234, B1 => n1992, B2 => 
                           n27230, ZN => n910_port);
   U1870 : OAI221_X1 port map( B1 => n1997, B2 => n27242, C1 => n1998, C2 => 
                           n27238, A => n892_port, ZN => n885_port);
   U1871 : AOI22_X1 port map( A1 => n1995, A2 => n27234, B1 => n1996, B2 => 
                           n27230, ZN => n892_port);
   U1872 : OAI221_X1 port map( B1 => n2001, B2 => n27242, C1 => n2002, C2 => 
                           n27238, A => n874_port, ZN => n867_port);
   U1873 : AOI22_X1 port map( A1 => n1999, A2 => n27234, B1 => n2000, B2 => 
                           n27230, ZN => n874_port);
   U1874 : OAI221_X1 port map( B1 => n2005, B2 => n27242, C1 => n2006, C2 => 
                           n27238, A => n856_port, ZN => n849_port);
   U1875 : AOI22_X1 port map( A1 => n2003, A2 => n27234, B1 => n2004, B2 => 
                           n27230, ZN => n856_port);
   U1876 : OAI221_X1 port map( B1 => n2009, B2 => n27243, C1 => n2010, C2 => 
                           n27239, A => n820_port, ZN => n813_port);
   U1877 : AOI22_X1 port map( A1 => n2007, A2 => n27234, B1 => n2008, B2 => 
                           n27230, ZN => n820_port);
   U1878 : OAI221_X1 port map( B1 => n2013, B2 => n27243, C1 => n2014, C2 => 
                           n27239, A => n798_port, ZN => n789_port);
   U1879 : AOI22_X1 port map( A1 => n2011, A2 => n27235, B1 => n2012, B2 => 
                           n27231, ZN => n798_port);
   U1880 : OAI221_X1 port map( B1 => n26359, B2 => n27139, C1 => n26632, C2 => 
                           n27135, A => n1862, ZN => n1847);
   U1881 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_0_port, B1 => n27127, 
                           B2 => regs_15_0_port, ZN => n1862);
   U1882 : OAI221_X1 port map( B1 => n26360, B2 => n27140, C1 => n26633, C2 => 
                           n27136, A => n1656, ZN => n1649);
   U1883 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_1_port, B1 => n27128, 
                           B2 => regs_15_1_port, ZN => n1656);
   U1884 : OAI221_X1 port map( B1 => n26361, B2 => n27141, C1 => n26634, C2 => 
                           n27137, A => n1458, ZN => n1451);
   U1885 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_2_port, B1 => n27129, 
                           B2 => regs_15_2_port, ZN => n1458);
   U1886 : OAI221_X1 port map( B1 => n26362, B2 => n27141, C1 => n26635, C2 => 
                           n27137, A => n1404, ZN => n1397);
   U1887 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_3_port, B1 => n27129, 
                           B2 => regs_15_3_port, ZN => n1404);
   U1888 : OAI221_X1 port map( B1 => n26363, B2 => n27141, C1 => n26636, C2 => 
                           n27137, A => n1386, ZN => n1379);
   U1889 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_4_port, B1 => n27129, 
                           B2 => regs_15_4_port, ZN => n1386);
   U1890 : OAI221_X1 port map( B1 => n26364, B2 => n27141, C1 => n26637, C2 => 
                           n27137, A => n1368, ZN => n1361);
   U1891 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_5_port, B1 => n27129, 
                           B2 => regs_15_5_port, ZN => n1368);
   U1892 : OAI221_X1 port map( B1 => n26365, B2 => n27141, C1 => n26638, C2 => 
                           n27137, A => n1350, ZN => n1343);
   U1893 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_6_port, B1 => n27129, 
                           B2 => regs_15_6_port, ZN => n1350);
   U1894 : OAI221_X1 port map( B1 => n26366, B2 => n27141, C1 => n26639, C2 => 
                           n27137, A => n1332, ZN => n1325);
   U1895 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_7_port, B1 => n27129, 
                           B2 => regs_15_7_port, ZN => n1332);
   U1896 : OAI221_X1 port map( B1 => n26367, B2 => n27141, C1 => n26640, C2 => 
                           n27137, A => n1314, ZN => n1307);
   U1897 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_8_port, B1 => n27129, 
                           B2 => regs_15_8_port, ZN => n1314);
   U1898 : OAI221_X1 port map( B1 => n26368, B2 => n27141, C1 => n26641, C2 => 
                           n27137, A => n1278, ZN => n1257);
   U1899 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_9_port, B1 => n27129, 
                           B2 => regs_15_9_port, ZN => n1278);
   U1900 : OAI221_X1 port map( B1 => n26369, B2 => n27139, C1 => n26642, C2 => 
                           n27135, A => n1836, ZN => n1829);
   U1901 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_10_port, B1 => n27127,
                           B2 => regs_15_10_port, ZN => n1836);
   U1902 : OAI221_X1 port map( B1 => n26370, B2 => n27139, C1 => n26643, C2 => 
                           n27135, A => n1818, ZN => n1811);
   U1903 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_11_port, B1 => n27127,
                           B2 => regs_15_11_port, ZN => n1818);
   U1904 : OAI221_X1 port map( B1 => n26371, B2 => n27139, C1 => n26644, C2 => 
                           n27135, A => n1800, ZN => n1793);
   U1905 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_12_port, B1 => n27127,
                           B2 => regs_15_12_port, ZN => n1800);
   U1906 : OAI221_X1 port map( B1 => n26372, B2 => n27139, C1 => n26645, C2 => 
                           n27135, A => n1782, ZN => n1775);
   U1907 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_13_port, B1 => n27127,
                           B2 => regs_15_13_port, ZN => n1782);
   U1908 : OAI221_X1 port map( B1 => n26373, B2 => n27139, C1 => n26646, C2 => 
                           n27135, A => n1764, ZN => n1757);
   U1909 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_14_port, B1 => n27127,
                           B2 => regs_15_14_port, ZN => n1764);
   U1910 : OAI221_X1 port map( B1 => n26374, B2 => n27139, C1 => n26647, C2 => 
                           n27135, A => n1746, ZN => n1739);
   U1911 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_15_port, B1 => n27127,
                           B2 => regs_15_15_port, ZN => n1746);
   U1912 : OAI221_X1 port map( B1 => n26375, B2 => n27139, C1 => n26648, C2 => 
                           n27135, A => n1728, ZN => n1721);
   U1913 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_16_port, B1 => n27127,
                           B2 => regs_15_16_port, ZN => n1728);
   U1914 : OAI221_X1 port map( B1 => n26376, B2 => n27139, C1 => n26649, C2 => 
                           n27135, A => n1710, ZN => n1703);
   U1915 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_17_port, B1 => n27127,
                           B2 => regs_15_17_port, ZN => n1710);
   U1916 : OAI221_X1 port map( B1 => n26377, B2 => n27139, C1 => n26650, C2 => 
                           n27135, A => n1692, ZN => n1685);
   U1917 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_18_port, B1 => n27127,
                           B2 => regs_15_18_port, ZN => n1692);
   U1918 : OAI221_X1 port map( B1 => n26378, B2 => n27139, C1 => n26651, C2 => 
                           n27135, A => n1674, ZN => n1667);
   U1919 : AOI22_X1 port map( A1 => n27131, A2 => regs_7_19_port, B1 => n27127,
                           B2 => regs_15_19_port, ZN => n1674);
   U1920 : OAI221_X1 port map( B1 => n26379, B2 => n27140, C1 => n26652, C2 => 
                           n27136, A => n1638, ZN => n1631);
   U1921 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_20_port, B1 => n27128,
                           B2 => regs_15_20_port, ZN => n1638);
   U1922 : OAI221_X1 port map( B1 => n26380, B2 => n27140, C1 => n26653, C2 => 
                           n27136, A => n1620, ZN => n1613);
   U1923 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_21_port, B1 => n27128,
                           B2 => regs_15_21_port, ZN => n1620);
   U1924 : OAI221_X1 port map( B1 => n26381, B2 => n27140, C1 => n26654, C2 => 
                           n27136, A => n1602, ZN => n1595);
   U1925 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_22_port, B1 => n27128,
                           B2 => regs_15_22_port, ZN => n1602);
   U1926 : OAI221_X1 port map( B1 => n26382, B2 => n27140, C1 => n26655, C2 => 
                           n27136, A => n1584, ZN => n1577);
   U1927 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_23_port, B1 => n27128,
                           B2 => regs_15_23_port, ZN => n1584);
   U1928 : OAI221_X1 port map( B1 => n26383, B2 => n27140, C1 => n26656, C2 => 
                           n27136, A => n1566, ZN => n1559);
   U1929 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_24_port, B1 => n27128,
                           B2 => regs_15_24_port, ZN => n1566);
   U1930 : OAI221_X1 port map( B1 => n26384, B2 => n27140, C1 => n26657, C2 => 
                           n27136, A => n1548, ZN => n1541);
   U1931 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_25_port, B1 => n27128,
                           B2 => regs_15_25_port, ZN => n1548);
   U1932 : OAI221_X1 port map( B1 => n26385, B2 => n27140, C1 => n26658, C2 => 
                           n27136, A => n1530, ZN => n1523);
   U1933 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_26_port, B1 => n27128,
                           B2 => regs_15_26_port, ZN => n1530);
   U1934 : OAI221_X1 port map( B1 => n26386, B2 => n27140, C1 => n26659, C2 => 
                           n27136, A => n1512, ZN => n1505);
   U1935 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_27_port, B1 => n27128,
                           B2 => regs_15_27_port, ZN => n1512);
   U1936 : OAI221_X1 port map( B1 => n26387, B2 => n27140, C1 => n26660, C2 => 
                           n27136, A => n1494, ZN => n1487);
   U1937 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_28_port, B1 => n27128,
                           B2 => regs_15_28_port, ZN => n1494);
   U1938 : OAI221_X1 port map( B1 => n26388, B2 => n27140, C1 => n26661, C2 => 
                           n27136, A => n1476, ZN => n1469);
   U1939 : AOI22_X1 port map( A1 => n27132, A2 => regs_7_29_port, B1 => n27128,
                           B2 => regs_15_29_port, ZN => n1476);
   U1940 : OAI221_X1 port map( B1 => n26389, B2 => n27141, C1 => n26662, C2 => 
                           n27137, A => n1440, ZN => n1433);
   U1941 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_30_port, B1 => n27129,
                           B2 => regs_15_30_port, ZN => n1440);
   U1942 : OAI221_X1 port map( B1 => n26390, B2 => n27141, C1 => n26663, C2 => 
                           n27137, A => n1422, ZN => n1415);
   U1943 : AOI22_X1 port map( A1 => n27133, A2 => regs_7_31_port, B1 => n27129,
                           B2 => regs_15_31_port, ZN => n1422);
   U1944 : AND2_X1 port map( A1 => add_rd2(3), A2 => add_rd2(4), ZN => n1232);
   U1945 : AOI22_X1 port map( A1 => n2639, A2 => n27705, B1 => n2638, B2 => 
                           n27706, ZN => n1254);
   U1946 : AOI22_X1 port map( A1 => n2641, A2 => n27705, B1 => n2640, B2 => 
                           n27706, ZN => n1044_port);
   U1947 : AOI22_X1 port map( A1 => n2643, A2 => n27705, B1 => n2642, B2 => 
                           n27706, ZN => n846_port);
   U1948 : AOI22_X1 port map( A1 => n2645, A2 => n27705, B1 => n2644, B2 => 
                           n27706, ZN => n786_port);
   U1949 : AOI22_X1 port map( A1 => n2647_port, A2 => n27705, B1 => n2646, B2 
                           => n27706, ZN => n768_port);
   U1950 : AOI22_X1 port map( A1 => n2288, A2 => n27705, B1 => n2287, B2 => 
                           n27706, ZN => n750_port);
   U1951 : AOI22_X1 port map( A1 => n2292, A2 => n27705, B1 => n2291, B2 => 
                           n27706, ZN => n732_port);
   U1952 : AOI22_X1 port map( A1 => n2296, A2 => n27705, B1 => n2295_port, B2 
                           => n27706, ZN => n714_port);
   U1953 : AOI22_X1 port map( A1 => n2300, A2 => n27705, B1 => n2299, B2 => 
                           n27706, ZN => n696_port);
   U1954 : AOI22_X1 port map( A1 => n2304, A2 => n27705, B1 => n2303, B2 => 
                           n27706, ZN => n678_port);
   U1955 : AOI22_X1 port map( A1 => n2308, A2 => n27705, B1 => n2307, B2 => 
                           n27706, ZN => n1224);
   U1956 : AOI22_X1 port map( A1 => n2312, A2 => n27705, B1 => n2311, B2 => 
                           n27706, ZN => n1206);
   U1957 : AOI22_X1 port map( A1 => n2316, A2 => n27705, B1 => n2315, B2 => 
                           n27706, ZN => n1188);
   U1958 : AOI22_X1 port map( A1 => n2320, A2 => n27705, B1 => n2319, B2 => 
                           n27706, ZN => n1170);
   U1959 : AOI22_X1 port map( A1 => n2324, A2 => n27705, B1 => n2323, B2 => 
                           n27706, ZN => n1152);
   U1960 : AOI22_X1 port map( A1 => n2328, A2 => n27705, B1 => n2327_port, B2 
                           => n27706, ZN => n1134);
   U1961 : AOI22_X1 port map( A1 => n2332, A2 => n27705, B1 => n2331, B2 => 
                           n27706, ZN => n1116);
   U1962 : AOI22_X1 port map( A1 => n2336, A2 => n27705, B1 => n2335, B2 => 
                           n27706, ZN => n1098);
   U1963 : AOI22_X1 port map( A1 => n2340, A2 => n27705, B1 => n2339, B2 => 
                           n27706, ZN => n1080);
   U1964 : AOI22_X1 port map( A1 => n2344, A2 => n27705, B1 => n2343, B2 => 
                           n27706, ZN => n1062);
   U1965 : AOI22_X1 port map( A1 => n2348, A2 => n27705, B1 => n2347, B2 => 
                           n27706, ZN => n1026_port);
   U1966 : AOI22_X1 port map( A1 => n2352, A2 => n27705, B1 => n2351, B2 => 
                           n27706, ZN => n1008_port);
   U1967 : AOI22_X1 port map( A1 => n2356, A2 => n27705, B1 => n2355, B2 => 
                           n27706, ZN => n990_port);
   U1968 : AOI22_X1 port map( A1 => regs_15_23_port, A2 => n27202, B1 => 
                           regs_7_23_port, B2 => n27198, ZN => n970_port);
   U1969 : AOI22_X1 port map( A1 => regs_15_24_port, A2 => n27202, B1 => 
                           regs_7_24_port, B2 => n27198, ZN => n952_port);
   U1970 : AOI22_X1 port map( A1 => regs_15_25_port, A2 => n27202, B1 => 
                           regs_7_25_port, B2 => n27198, ZN => n934_port);
   U1971 : AOI22_X1 port map( A1 => regs_15_26_port, A2 => n27202, B1 => 
                           regs_7_26_port, B2 => n27198, ZN => n916_port);
   U1972 : AOI22_X1 port map( A1 => regs_15_27_port, A2 => n27202, B1 => 
                           regs_7_27_port, B2 => n27198, ZN => n898_port);
   U1973 : AOI22_X1 port map( A1 => regs_15_28_port, A2 => n27202, B1 => 
                           regs_7_28_port, B2 => n27198, ZN => n880_port);
   U1974 : AOI22_X1 port map( A1 => regs_15_29_port, A2 => n27202, B1 => 
                           regs_7_29_port, B2 => n27198, ZN => n862_port);
   U1975 : AOI22_X1 port map( A1 => regs_15_30_port, A2 => n27202, B1 => 
                           regs_7_30_port, B2 => n27198, ZN => n826_port);
   U1976 : AOI22_X1 port map( A1 => regs_15_31_port, A2 => n27203, B1 => 
                           regs_7_31_port, B2 => n27199, ZN => n804_port);
   U1977 : AOI22_X1 port map( A1 => n27067, A2 => n26443, B1 => n27063, B2 => 
                           n26782, ZN => n1874);
   U1978 : AOI22_X1 port map( A1 => n27068, A2 => n26444, B1 => n27064, B2 => 
                           n26783, ZN => n1664);
   U1979 : AOI22_X1 port map( A1 => n27069, A2 => n26445, B1 => n27065, B2 => 
                           n26784, ZN => n1466);
   U1980 : AOI22_X1 port map( A1 => n27069, A2 => n26446, B1 => n27065, B2 => 
                           n26785, ZN => n1412);
   U1981 : AOI22_X1 port map( A1 => n27069, A2 => n26447, B1 => n27065, B2 => 
                           n26786, ZN => n1394);
   U1982 : AOI22_X1 port map( A1 => n27069, A2 => n26448, B1 => n27065, B2 => 
                           n26787, ZN => n1376);
   U1983 : AOI22_X1 port map( A1 => n27069, A2 => n26449, B1 => n27065, B2 => 
                           n26788, ZN => n1358);
   U1984 : AOI22_X1 port map( A1 => n27069, A2 => n26450, B1 => n27065, B2 => 
                           n26789, ZN => n1340);
   U1985 : AOI22_X1 port map( A1 => n27069, A2 => n26451, B1 => n27065, B2 => 
                           n26790, ZN => n1322);
   U1986 : AOI22_X1 port map( A1 => n27069, A2 => n26452, B1 => n27065, B2 => 
                           n26791, ZN => n1302);
   U1987 : AOI22_X1 port map( A1 => n27067, A2 => n26453, B1 => n27063, B2 => 
                           n26792, ZN => n1844);
   U1988 : AOI22_X1 port map( A1 => n27067, A2 => n26454, B1 => n27063, B2 => 
                           n26793, ZN => n1826);
   U1989 : AOI22_X1 port map( A1 => n27067, A2 => n26455, B1 => n27063, B2 => 
                           n26794, ZN => n1808);
   U1990 : AOI22_X1 port map( A1 => n27067, A2 => n26456, B1 => n27063, B2 => 
                           n26795, ZN => n1790);
   U1991 : AOI22_X1 port map( A1 => n27067, A2 => n26457, B1 => n27063, B2 => 
                           n26796, ZN => n1772);
   U1992 : AOI22_X1 port map( A1 => n27067, A2 => n26458, B1 => n27063, B2 => 
                           n26797, ZN => n1754);
   U1993 : AOI22_X1 port map( A1 => n27067, A2 => n26459, B1 => n27063, B2 => 
                           n26798, ZN => n1736);
   U1994 : AOI22_X1 port map( A1 => n27067, A2 => n26460, B1 => n27063, B2 => 
                           n26799, ZN => n1718);
   U1995 : AOI22_X1 port map( A1 => n27067, A2 => n26461, B1 => n27063, B2 => 
                           n26800, ZN => n1700);
   U1996 : AOI22_X1 port map( A1 => n27067, A2 => n26462, B1 => n27063, B2 => 
                           n26801, ZN => n1682);
   U1997 : AOI22_X1 port map( A1 => n27068, A2 => n26463, B1 => n27064, B2 => 
                           n26802, ZN => n1646);
   U1998 : AOI22_X1 port map( A1 => n27068, A2 => n26464, B1 => n27064, B2 => 
                           n26803, ZN => n1628);
   U1999 : AOI22_X1 port map( A1 => n27068, A2 => n26465, B1 => n27064, B2 => 
                           n26804, ZN => n1610);
   U2000 : AOI22_X1 port map( A1 => n27068, A2 => n26466, B1 => n27064, B2 => 
                           n26805, ZN => n1592);
   U2001 : AOI22_X1 port map( A1 => n27068, A2 => n26467, B1 => n27064, B2 => 
                           n26806, ZN => n1574);
   U2002 : AOI22_X1 port map( A1 => n27068, A2 => n26468, B1 => n27064, B2 => 
                           n26807, ZN => n1556);
   U2003 : AOI22_X1 port map( A1 => n27068, A2 => n26469, B1 => n27064, B2 => 
                           n26808, ZN => n1538);
   U2004 : AOI22_X1 port map( A1 => n27068, A2 => n26470, B1 => n27064, B2 => 
                           n26809, ZN => n1520);
   U2005 : AOI22_X1 port map( A1 => n27068, A2 => n26471, B1 => n27064, B2 => 
                           n26810, ZN => n1502);
   U2006 : AOI22_X1 port map( A1 => n27068, A2 => n26472, B1 => n27064, B2 => 
                           n26811, ZN => n1484);
   U2007 : AOI22_X1 port map( A1 => n27069, A2 => n26473, B1 => n27065, B2 => 
                           n26812, ZN => n1448);
   U2008 : AOI22_X1 port map( A1 => n27069, A2 => n26474, B1 => n27065, B2 => 
                           n26813, ZN => n1430);
   U2009 : INV_X1 port map( A => add_rd1(2), ZN => n27717);
   U2010 : INV_X1 port map( A => add_rd2(2), ZN => n27713);
   U2011 : INV_X1 port map( A => add_rd1(1), ZN => n27716);
   U2012 : INV_X1 port map( A => add_rd2(1), ZN => n27712);
   U2013 : INV_X1 port map( A => add_rd1(0), ZN => n27715);
   U2014 : INV_X1 port map( A => add_rd2(0), ZN => n27704);
   U2015 : INV_X1 port map( A => add_wr(2), ZN => n27698);
   U2016 : INV_X1 port map( A => add_wr(0), ZN => n27696);
   U2017 : INV_X1 port map( A => add_wr(1), ZN => n27697);
   U2018 : INV_X1 port map( A => n1196, ZN => n27695);
   U2019 : AOI221_X1 port map( B1 => n27703, B2 => n25445, C1 => n26589, C2 => 
                           n27702, A => n1197, ZN => n1196);
   U2020 : OAI22_X1 port map( A1 => n651_port, A2 => n25511, B1 => n26596, B2 
                           => n652_port, ZN => n1197);
   U2021 : INV_X1 port map( A => n1178, ZN => n27694);
   U2022 : AOI221_X1 port map( B1 => n27703, B2 => n25446, C1 => n26590, C2 => 
                           n27702, A => n1179, ZN => n1178);
   U2023 : OAI22_X1 port map( A1 => n651_port, A2 => n25512, B1 => n26597, B2 
                           => n652_port, ZN => n1179);
   U2024 : INV_X1 port map( A => n1160, ZN => n27693);
   U2025 : AOI221_X1 port map( B1 => n27703, B2 => n25447, C1 => n26591, C2 => 
                           n27702, A => n1161, ZN => n1160);
   U2026 : OAI22_X1 port map( A1 => n651_port, A2 => n25513, B1 => n26598, B2 
                           => n652_port, ZN => n1161);
   U2027 : INV_X1 port map( A => n1142, ZN => n27692);
   U2028 : AOI221_X1 port map( B1 => n27703, B2 => n25448, C1 => n26592, C2 => 
                           n27702, A => n1143, ZN => n1142);
   U2029 : OAI22_X1 port map( A1 => n651_port, A2 => n25514, B1 => n26599, B2 
                           => n652_port, ZN => n1143);
   U2030 : INV_X1 port map( A => add_rd1(3), ZN => n27718);
   U2031 : INV_X1 port map( A => add_rd1(4), ZN => n27719);
   U2032 : NAND2_X1 port map( A1 => n1009_port, A2 => n1010_port, ZN => 
                           out2(20));
   U2033 : NOR4_X1 port map( A1 => n1019_port, A2 => n1020_port, A3 => 
                           n1021_port, A4 => n1022_port, ZN => n1009_port);
   U2034 : NOR4_X1 port map( A1 => n1011_port, A2 => n1012_port, A3 => 
                           n1013_port, A4 => n1014_port, ZN => n1010_port);
   U2035 : OAI221_X1 port map( B1 => n2349, B2 => n27193, C1 => n2350, C2 => 
                           n27190, A => n1026_port, ZN => n1019_port);
   U2036 : NAND2_X1 port map( A1 => n991_port, A2 => n992_port, ZN => out2(21))
                           ;
   U2037 : NOR4_X1 port map( A1 => n1001_port, A2 => n1002_port, A3 => 
                           n1003_port, A4 => n1004_port, ZN => n991_port);
   U2038 : NOR4_X1 port map( A1 => n993_port, A2 => n994_port, A3 => n995_port,
                           A4 => n996_port, ZN => n992_port);
   U2039 : OAI221_X1 port map( B1 => n2353, B2 => n27193, C1 => n2354, C2 => 
                           n27190, A => n1008_port, ZN => n1001_port);
   U2040 : NAND2_X1 port map( A1 => n973_port, A2 => n974_port, ZN => out2(22))
                           ;
   U2041 : NOR4_X1 port map( A1 => n983_port, A2 => n984_port, A3 => n985_port,
                           A4 => n986_port, ZN => n973_port);
   U2042 : NOR4_X1 port map( A1 => n975_port, A2 => n976_port, A3 => n977_port,
                           A4 => n978_port, ZN => n974_port);
   U2043 : OAI221_X1 port map( B1 => n2357, B2 => n27193, C1 => n2358, C2 => 
                           n27190, A => n990_port, ZN => n983_port);
   U2044 : NAND2_X1 port map( A1 => n1225, A2 => n1226, ZN => out2(0));
   U2045 : NOR4_X1 port map( A1 => n1245, A2 => n1246, A3 => n1247, A4 => n1248
                           , ZN => n1225);
   U2046 : NOR4_X1 port map( A1 => n1227, A2 => n1228, A3 => n1229, A4 => n1230
                           , ZN => n1226);
   U2047 : OAI221_X1 port map( B1 => n2649, B2 => n27193, C1 => n2648, C2 => 
                           n27190, A => n1254, ZN => n1245);
   U2048 : NAND2_X1 port map( A1 => n1027_port, A2 => n1028_port, ZN => out2(1)
                           );
   U2049 : NOR4_X1 port map( A1 => n1037_port, A2 => n1038_port, A3 => 
                           n1039_port, A4 => n1040_port, ZN => n1027_port);
   U2050 : NOR4_X1 port map( A1 => n1029_port, A2 => n1030_port, A3 => 
                           n1031_port, A4 => n1032_port, ZN => n1028_port);
   U2051 : OAI221_X1 port map( B1 => n2651, B2 => n27193, C1 => n2650, C2 => 
                           n27190, A => n1044_port, ZN => n1037_port);
   U2052 : NAND2_X1 port map( A1 => n829_port, A2 => n830_port, ZN => out2(2));
   U2053 : NOR4_X1 port map( A1 => n839_port, A2 => n840_port, A3 => n841_port,
                           A4 => n842_port, ZN => n829_port);
   U2054 : NOR4_X1 port map( A1 => n831_port, A2 => n832_port, A3 => n833_port,
                           A4 => n834_port, ZN => n830_port);
   U2055 : OAI221_X1 port map( B1 => n2653, B2 => n27193, C1 => n2652, C2 => 
                           n27190, A => n846_port, ZN => n839_port);
   U2056 : NAND2_X1 port map( A1 => n769_port, A2 => n770_port, ZN => out2(3));
   U2057 : NOR4_X1 port map( A1 => n779_port, A2 => n780_port, A3 => n781_port,
                           A4 => n782_port, ZN => n769_port);
   U2058 : NOR4_X1 port map( A1 => n771_port, A2 => n772_port, A3 => n773_port,
                           A4 => n774_port, ZN => n770_port);
   U2059 : OAI221_X1 port map( B1 => n2655, B2 => n27193, C1 => n2654, C2 => 
                           n27190, A => n786_port, ZN => n779_port);
   U2060 : NAND2_X1 port map( A1 => n751_port, A2 => n752_port, ZN => out2(4));
   U2061 : NOR4_X1 port map( A1 => n761_port, A2 => n762_port, A3 => n763_port,
                           A4 => n764_port, ZN => n751_port);
   U2062 : NOR4_X1 port map( A1 => n753_port, A2 => n754_port, A3 => n755_port,
                           A4 => n756_port, ZN => n752_port);
   U2063 : OAI221_X1 port map( B1 => n2657, B2 => n27193, C1 => n2656, C2 => 
                           n27190, A => n768_port, ZN => n761_port);
   U2064 : NAND2_X1 port map( A1 => n733_port, A2 => n734_port, ZN => out2(5));
   U2065 : NOR4_X1 port map( A1 => n743_port, A2 => n744_port, A3 => n745_port,
                           A4 => n746_port, ZN => n733_port);
   U2066 : NOR4_X1 port map( A1 => n735_port, A2 => n736_port, A3 => n737_port,
                           A4 => n738_port, ZN => n734_port);
   U2067 : OAI221_X1 port map( B1 => n2289, B2 => n27193, C1 => n2290, C2 => 
                           n27190, A => n750_port, ZN => n743_port);
   U2068 : NAND2_X1 port map( A1 => n715_port, A2 => n716_port, ZN => out2(6));
   U2069 : NOR4_X1 port map( A1 => n725_port, A2 => n726_port, A3 => n727_port,
                           A4 => n728_port, ZN => n715_port);
   U2070 : NOR4_X1 port map( A1 => n717_port, A2 => n718_port, A3 => n719_port,
                           A4 => n720_port, ZN => n716_port);
   U2071 : OAI221_X1 port map( B1 => n2293, B2 => n27193, C1 => n2294, C2 => 
                           n27190, A => n732_port, ZN => n725_port);
   U2072 : NAND2_X1 port map( A1 => n697_port, A2 => n698_port, ZN => out2(7));
   U2073 : NOR4_X1 port map( A1 => n707_port, A2 => n708_port, A3 => n709_port,
                           A4 => n710_port, ZN => n697_port);
   U2074 : NOR4_X1 port map( A1 => n699_port, A2 => n700_port, A3 => n701_port,
                           A4 => n702_port, ZN => n698_port);
   U2075 : OAI221_X1 port map( B1 => n2297, B2 => n27193, C1 => n2298, C2 => 
                           n27190, A => n714_port, ZN => n707_port);
   U2076 : NAND2_X1 port map( A1 => n679_port, A2 => n680_port, ZN => out2(8));
   U2077 : NOR4_X1 port map( A1 => n689_port, A2 => n690_port, A3 => n691_port,
                           A4 => n692_port, ZN => n679_port);
   U2078 : NOR4_X1 port map( A1 => n681_port, A2 => n682_port, A3 => n683_port,
                           A4 => n684_port, ZN => n680_port);
   U2079 : OAI221_X1 port map( B1 => n2301, B2 => n27193, C1 => n2302, C2 => 
                           n27190, A => n696_port, ZN => n689_port);
   U2080 : NAND2_X1 port map( A1 => n635_port, A2 => n636_port, ZN => out2(9));
   U2081 : NOR4_X1 port map( A1 => n659_port, A2 => n660_port, A3 => n661_port,
                           A4 => n662_port, ZN => n635_port);
   U2082 : NOR4_X1 port map( A1 => n637_port, A2 => n638_port, A3 => n639_port,
                           A4 => n640_port, ZN => n636_port);
   U2083 : OAI221_X1 port map( B1 => n2305, B2 => n27193, C1 => n2306, C2 => 
                           n27190, A => n678_port, ZN => n659_port);
   U2084 : NAND2_X1 port map( A1 => n1207, A2 => n1208, ZN => out2(10));
   U2085 : NOR4_X1 port map( A1 => n1217, A2 => n1218, A3 => n1219, A4 => n1220
                           , ZN => n1207);
   U2086 : NOR4_X1 port map( A1 => n1209, A2 => n1210, A3 => n1211, A4 => n1212
                           , ZN => n1208);
   U2087 : OAI221_X1 port map( B1 => n2309, B2 => n27193, C1 => n2310, C2 => 
                           n27190, A => n1224, ZN => n1217);
   U2088 : NAND2_X1 port map( A1 => n1189, A2 => n1190, ZN => out2(11));
   U2089 : NOR4_X1 port map( A1 => n1199, A2 => n1200, A3 => n1201, A4 => n1202
                           , ZN => n1189);
   U2090 : NOR4_X1 port map( A1 => n1191, A2 => n27695, A3 => n1192, A4 => 
                           n1193, ZN => n1190);
   U2091 : OAI221_X1 port map( B1 => n2313, B2 => n27193, C1 => n2314, C2 => 
                           n27190, A => n1206, ZN => n1199);
   U2092 : NAND2_X1 port map( A1 => n1171, A2 => n1172, ZN => out2(12));
   U2093 : NOR4_X1 port map( A1 => n1181, A2 => n1182, A3 => n1183, A4 => n1184
                           , ZN => n1171);
   U2094 : NOR4_X1 port map( A1 => n1173, A2 => n27694, A3 => n1174, A4 => 
                           n1175, ZN => n1172);
   U2095 : OAI221_X1 port map( B1 => n2317, B2 => n27193, C1 => n2318, C2 => 
                           n27190, A => n1188, ZN => n1181);
   U2096 : NAND2_X1 port map( A1 => n1153, A2 => n1154, ZN => out2(13));
   U2097 : NOR4_X1 port map( A1 => n1163, A2 => n1164, A3 => n1165, A4 => n1166
                           , ZN => n1153);
   U2098 : NOR4_X1 port map( A1 => n1155, A2 => n27693, A3 => n1156, A4 => 
                           n1157, ZN => n1154);
   U2099 : OAI221_X1 port map( B1 => n2321, B2 => n27193, C1 => n2322, C2 => 
                           n27190, A => n1170, ZN => n1163);
   U2100 : NAND2_X1 port map( A1 => n1135, A2 => n1136, ZN => out2(14));
   U2101 : NOR4_X1 port map( A1 => n1145, A2 => n1146, A3 => n1147, A4 => n1148
                           , ZN => n1135);
   U2102 : NOR4_X1 port map( A1 => n1137, A2 => n27692, A3 => n1138, A4 => 
                           n1139, ZN => n1136);
   U2103 : OAI221_X1 port map( B1 => n2325, B2 => n27193, C1 => n2326, C2 => 
                           n27190, A => n1152, ZN => n1145);
   U2104 : NAND2_X1 port map( A1 => n1117, A2 => n1118, ZN => out2(15));
   U2105 : NOR4_X1 port map( A1 => n1127, A2 => n1128, A3 => n1129, A4 => n1130
                           , ZN => n1117);
   U2106 : NOR4_X1 port map( A1 => n1119, A2 => n1120, A3 => n1121, A4 => n1122
                           , ZN => n1118);
   U2107 : OAI221_X1 port map( B1 => n2329, B2 => n27193, C1 => n2330, C2 => 
                           n27190, A => n1134, ZN => n1127);
   U2108 : NAND2_X1 port map( A1 => n1099, A2 => n1100, ZN => out2(16));
   U2109 : NOR4_X1 port map( A1 => n1109, A2 => n1110, A3 => n1111, A4 => n1112
                           , ZN => n1099);
   U2110 : NOR4_X1 port map( A1 => n1101, A2 => n1102, A3 => n1103, A4 => n1104
                           , ZN => n1100);
   U2111 : OAI221_X1 port map( B1 => n2333, B2 => n27193, C1 => n2334, C2 => 
                           n27190, A => n1116, ZN => n1109);
   U2112 : NAND2_X1 port map( A1 => n1081, A2 => n1082, ZN => out2(17));
   U2113 : NOR4_X1 port map( A1 => n1091, A2 => n1092, A3 => n1093, A4 => n1094
                           , ZN => n1081);
   U2114 : NOR4_X1 port map( A1 => n1083, A2 => n1084, A3 => n1085, A4 => n1086
                           , ZN => n1082);
   U2115 : OAI221_X1 port map( B1 => n2337, B2 => n27193, C1 => n2338, C2 => 
                           n27190, A => n1098, ZN => n1091);
   U2116 : NAND2_X1 port map( A1 => n1063, A2 => n1064, ZN => out2(18));
   U2117 : NOR4_X1 port map( A1 => n1073, A2 => n1074, A3 => n1075, A4 => n1076
                           , ZN => n1063);
   U2118 : NOR4_X1 port map( A1 => n1065, A2 => n1066, A3 => n1067, A4 => n1068
                           , ZN => n1064);
   U2119 : OAI221_X1 port map( B1 => n2341, B2 => n27193, C1 => n2342, C2 => 
                           n27190, A => n1080, ZN => n1073);
   U2120 : NAND2_X1 port map( A1 => n1045_port, A2 => n1046_port, ZN => 
                           out2(19));
   U2121 : NOR4_X1 port map( A1 => n1055, A2 => n1056, A3 => n1057, A4 => n1058
                           , ZN => n1045_port);
   U2122 : NOR4_X1 port map( A1 => n1047, A2 => n1048, A3 => n1049, A4 => n1050
                           , ZN => n1046_port);
   U2123 : OAI221_X1 port map( B1 => n2345, B2 => n27193, C1 => n2346, C2 => 
                           n27190, A => n1062, ZN => n1055);
   U2124 : INV_X1 port map( A => add_rd2(3), ZN => n27714);
   U2125 : INV_X1 port map( A => rst, ZN => n27720);
   U2126 : INV_X1 port map( A => add_wr(4), ZN => n27700);
   U2127 : INV_X1 port map( A => add_wr(3), ZN => n27699);
   U2128 : AND2_X1 port map( A1 => regs_nxt_31_0_port, A2 => n27006, ZN => N23)
                           ;
   U2129 : AND2_X1 port map( A1 => regs_nxt_31_1_port, A2 => n27007, ZN => N24)
                           ;
   U2130 : AND2_X1 port map( A1 => regs_nxt_31_2_port, A2 => n27007, ZN => N25)
                           ;
   U2131 : AND2_X1 port map( A1 => regs_nxt_31_3_port, A2 => n27008, ZN => N26)
                           ;
   U2132 : AND2_X1 port map( A1 => regs_nxt_31_4_port, A2 => n27009, ZN => N27)
                           ;
   U2133 : AND2_X1 port map( A1 => regs_nxt_31_5_port, A2 => n27009, ZN => N28)
                           ;
   U2134 : AND2_X1 port map( A1 => regs_nxt_31_6_port, A2 => n27010, ZN => N29)
                           ;
   U2135 : AND2_X1 port map( A1 => regs_nxt_31_7_port, A2 => n27011, ZN => N30)
                           ;
   U2136 : AND2_X1 port map( A1 => regs_nxt_31_8_port, A2 => n27029, ZN => N31)
                           ;
   U2137 : AND2_X1 port map( A1 => regs_nxt_31_9_port, A2 => n27026, ZN => N32)
                           ;
   U2138 : AND2_X1 port map( A1 => regs_nxt_31_10_port, A2 => n27027, ZN => N33
                           );
   U2139 : AND2_X1 port map( A1 => regs_nxt_31_11_port, A2 => n27028, ZN => N34
                           );
   U2140 : AND2_X1 port map( A1 => regs_nxt_31_12_port, A2 => n27028, ZN => N35
                           );
   U2141 : AND2_X1 port map( A1 => regs_nxt_31_13_port, A2 => n27029, ZN => N36
                           );
   U2142 : AND2_X1 port map( A1 => regs_nxt_31_14_port, A2 => n27029, ZN => N37
                           );
   U2143 : AND2_X1 port map( A1 => regs_nxt_31_15_port, A2 => n27030, ZN => N38
                           );
   U2144 : AND2_X1 port map( A1 => regs_nxt_31_16_port, A2 => n27031, ZN => N39
                           );
   U2145 : AND2_X1 port map( A1 => regs_nxt_31_17_port, A2 => n27031, ZN => N40
                           );
   U2146 : AND2_X1 port map( A1 => regs_nxt_31_18_port, A2 => n27032, ZN => N41
                           );
   U2147 : AND2_X1 port map( A1 => regs_nxt_31_19_port, A2 => n27033, ZN => N42
                           );
   U2148 : AND2_X1 port map( A1 => regs_nxt_31_20_port, A2 => n27018, ZN => N43
                           );
   U2149 : AND2_X1 port map( A1 => regs_nxt_31_21_port, A2 => n27019, ZN => N44
                           );
   U2150 : AND2_X1 port map( A1 => regs_nxt_31_22_port, A2 => n27020, ZN => N45
                           );
   U2151 : AND2_X1 port map( A1 => regs_nxt_31_23_port, A2 => n27020, ZN => N46
                           );
   U2152 : AND2_X1 port map( A1 => regs_nxt_31_24_port, A2 => n27021, ZN => N47
                           );
   U2153 : AND2_X1 port map( A1 => regs_nxt_31_25_port, A2 => n27022, ZN => N48
                           );
   U2154 : AND2_X1 port map( A1 => regs_nxt_31_26_port, A2 => n27022, ZN => N49
                           );
   U2155 : AND2_X1 port map( A1 => regs_nxt_31_27_port, A2 => n27023, ZN => N50
                           );
   U2156 : AND2_X1 port map( A1 => regs_nxt_31_28_port, A2 => n27023, ZN => N51
                           );
   U2157 : AND2_X1 port map( A1 => regs_nxt_31_29_port, A2 => n27024, ZN => N52
                           );
   U2158 : AND2_X1 port map( A1 => regs_nxt_31_30_port, A2 => n27025, ZN => N53
                           );
   U2159 : AND2_X1 port map( A1 => regs_nxt_31_31_port, A2 => n27025, ZN => N54
                           );
   U2160 : AND2_X1 port map( A1 => regs_nxt_30_0_port, A2 => n26974, ZN => N55)
                           ;
   U2161 : AND2_X1 port map( A1 => regs_nxt_30_1_port, A2 => n26981, ZN => N56)
                           ;
   U2162 : AND2_X1 port map( A1 => regs_nxt_30_2_port, A2 => n26982, ZN => N57)
                           ;
   U2163 : AND2_X1 port map( A1 => regs_nxt_30_3_port, A2 => n26983, ZN => N58)
                           ;
   U2164 : AND2_X1 port map( A1 => regs_nxt_30_4_port, A2 => n26983, ZN => N59)
                           ;
   U2165 : AND2_X1 port map( A1 => regs_nxt_30_5_port, A2 => n26984, ZN => N60)
                           ;
   U2166 : AND2_X1 port map( A1 => regs_nxt_30_6_port, A2 => n26984, ZN => N61)
                           ;
   U2167 : AND2_X1 port map( A1 => regs_nxt_30_7_port, A2 => n26985, ZN => N62)
                           ;
   U2168 : AND2_X1 port map( A1 => regs_nxt_30_8_port, A2 => n26986, ZN => N63)
                           ;
   U2169 : AND2_X1 port map( A1 => regs_nxt_30_9_port, A2 => n26986, ZN => N64)
                           ;
   U2170 : AND2_X1 port map( A1 => regs_nxt_30_10_port, A2 => n26987, ZN => N65
                           );
   U2171 : AND2_X1 port map( A1 => regs_nxt_30_11_port, A2 => n26988, ZN => N66
                           );
   U2172 : AND2_X1 port map( A1 => regs_nxt_30_12_port, A2 => n26988, ZN => N67
                           );
   U2173 : AND2_X1 port map( A1 => regs_nxt_30_13_port, A2 => n26989, ZN => N68
                           );
   U2174 : AND2_X1 port map( A1 => regs_nxt_30_14_port, A2 => n26975, ZN => N69
                           );
   U2175 : AND2_X1 port map( A1 => regs_nxt_30_15_port, A2 => n26975, ZN => N70
                           );
   U2176 : AND2_X1 port map( A1 => regs_nxt_30_16_port, A2 => n26976, ZN => N71
                           );
   U2177 : AND2_X1 port map( A1 => regs_nxt_30_17_port, A2 => n26977, ZN => N72
                           );
   U2178 : AND2_X1 port map( A1 => regs_nxt_30_18_port, A2 => n26977, ZN => N73
                           );
   U2179 : AND2_X1 port map( A1 => regs_nxt_30_19_port, A2 => n26978, ZN => N74
                           );
   U2180 : AND2_X1 port map( A1 => regs_nxt_30_20_port, A2 => n26979, ZN => N75
                           );
   U2181 : AND2_X1 port map( A1 => regs_nxt_30_21_port, A2 => n26979, ZN => N76
                           );
   U2182 : AND2_X1 port map( A1 => regs_nxt_30_22_port, A2 => n26980, ZN => N77
                           );
   U2183 : AND2_X1 port map( A1 => regs_nxt_30_23_port, A2 => n26980, ZN => N78
                           );
   U2184 : AND2_X1 port map( A1 => regs_nxt_30_24_port, A2 => n26996, ZN => N79
                           );
   U2185 : AND2_X1 port map( A1 => regs_nxt_30_25_port, A2 => n26997, ZN => N80
                           );
   U2186 : AND2_X1 port map( A1 => regs_nxt_30_26_port, A2 => n26998, ZN => N81
                           );
   U2187 : AND2_X1 port map( A1 => regs_nxt_30_27_port, A2 => n26998, ZN => N82
                           );
   U2188 : AND2_X1 port map( A1 => regs_nxt_30_28_port, A2 => n26999, ZN => N83
                           );
   U2189 : AND2_X1 port map( A1 => regs_nxt_30_29_port, A2 => n27000, ZN => N84
                           );
   U2190 : AND2_X1 port map( A1 => regs_nxt_30_30_port, A2 => n27000, ZN => N85
                           );
   U2191 : AND2_X1 port map( A1 => regs_nxt_30_31_port, A2 => n27001, ZN => N86
                           );
   U2192 : AND2_X1 port map( A1 => regs_nxt_29_0_port, A2 => n27001, ZN => N87)
                           ;
   U2193 : AND2_X1 port map( A1 => regs_nxt_29_1_port, A2 => n27002, ZN => N88)
                           ;
   U2194 : AND2_X1 port map( A1 => regs_nxt_29_2_port, A2 => n27003, ZN => N89)
                           ;
   U2195 : AND2_X1 port map( A1 => regs_nxt_29_3_port, A2 => n27003, ZN => N90)
                           ;
   U2196 : AND2_X1 port map( A1 => regs_nxt_29_4_port, A2 => n26989, ZN => N91)
                           ;
   U2197 : AND2_X1 port map( A1 => regs_nxt_29_5_port, A2 => n26990, ZN => N92)
                           ;
   U2198 : AND2_X1 port map( A1 => regs_nxt_29_6_port, A2 => n26990, ZN => N93)
                           ;
   U2199 : AND2_X1 port map( A1 => regs_nxt_29_7_port, A2 => n26991, ZN => N94)
                           ;
   U2200 : AND2_X1 port map( A1 => regs_nxt_29_8_port, A2 => n26992, ZN => N95)
                           ;
   U2201 : AND2_X1 port map( A1 => regs_nxt_29_9_port, A2 => n26992, ZN => N96)
                           ;
   U2202 : AND2_X1 port map( A1 => regs_nxt_29_10_port, A2 => n26993, ZN => N97
                           );
   U2203 : AND2_X1 port map( A1 => regs_nxt_29_11_port, A2 => n26993, ZN => N98
                           );
   U2204 : AND2_X1 port map( A1 => regs_nxt_29_12_port, A2 => n26994, ZN => N99
                           );
   U2205 : AND2_X1 port map( A1 => regs_nxt_29_13_port, A2 => n26981, ZN => 
                           N100);
   U2206 : AND2_X1 port map( A1 => regs_nxt_29_14_port, A2 => n27012, ZN => 
                           N101);
   U2207 : AND2_X1 port map( A1 => regs_nxt_29_15_port, A2 => n27012, ZN => 
                           N102);
   U2208 : AND2_X1 port map( A1 => regs_nxt_29_16_port, A2 => n27013, ZN => 
                           N103);
   U2209 : AND2_X1 port map( A1 => regs_nxt_29_17_port, A2 => n27013, ZN => 
                           N104);
   U2210 : AND2_X1 port map( A1 => regs_nxt_29_18_port, A2 => n27014, ZN => 
                           N105);
   U2211 : AND2_X1 port map( A1 => regs_nxt_29_19_port, A2 => n27014, ZN => 
                           N106);
   U2212 : AND2_X1 port map( A1 => regs_nxt_29_20_port, A2 => n27014, ZN => 
                           N107);
   U2213 : AND2_X1 port map( A1 => regs_nxt_29_21_port, A2 => n27014, ZN => 
                           N108);
   U2214 : AND2_X1 port map( A1 => regs_nxt_29_22_port, A2 => n27014, ZN => 
                           N109);
   U2215 : AND2_X1 port map( A1 => regs_nxt_29_23_port, A2 => n27014, ZN => 
                           N110);
   U2216 : AND2_X1 port map( A1 => regs_nxt_29_24_port, A2 => n27014, ZN => 
                           N111);
   U2217 : AND2_X1 port map( A1 => regs_nxt_29_25_port, A2 => n27014, ZN => 
                           N112);
   U2218 : AND2_X1 port map( A1 => regs_nxt_29_26_port, A2 => n27014, ZN => 
                           N113);
   U2219 : AND2_X1 port map( A1 => regs_nxt_29_27_port, A2 => n27014, ZN => 
                           N114);
   U2220 : AND2_X1 port map( A1 => regs_nxt_29_28_port, A2 => n27014, ZN => 
                           N115);
   U2221 : AND2_X1 port map( A1 => regs_nxt_29_29_port, A2 => n27014, ZN => 
                           N116);
   U2222 : AND2_X1 port map( A1 => regs_nxt_29_30_port, A2 => n27015, ZN => 
                           N117);
   U2223 : AND2_X1 port map( A1 => regs_nxt_29_31_port, A2 => n27015, ZN => 
                           N118);
   U2224 : AND2_X1 port map( A1 => regs_nxt_28_0_port, A2 => n27015, ZN => N119
                           );
   U2225 : AND2_X1 port map( A1 => regs_nxt_28_1_port, A2 => n27015, ZN => N120
                           );
   U2226 : AND2_X1 port map( A1 => regs_nxt_28_2_port, A2 => n27015, ZN => N121
                           );
   U2227 : AND2_X1 port map( A1 => regs_nxt_28_3_port, A2 => n27015, ZN => N122
                           );
   U2228 : AND2_X1 port map( A1 => regs_nxt_28_4_port, A2 => n27015, ZN => N123
                           );
   U2229 : AND2_X1 port map( A1 => regs_nxt_28_5_port, A2 => n27015, ZN => N124
                           );
   U2230 : AND2_X1 port map( A1 => regs_nxt_28_6_port, A2 => n27015, ZN => N125
                           );
   U2231 : AND2_X1 port map( A1 => regs_nxt_28_7_port, A2 => n27015, ZN => N126
                           );
   U2232 : AND2_X1 port map( A1 => regs_nxt_28_8_port, A2 => n27015, ZN => N127
                           );
   U2233 : AND2_X1 port map( A1 => regs_nxt_28_9_port, A2 => n27015, ZN => N128
                           );
   U2234 : AND2_X1 port map( A1 => regs_nxt_28_10_port, A2 => n27015, ZN => 
                           N129);
   U2235 : AND2_X1 port map( A1 => regs_nxt_28_11_port, A2 => n27015, ZN => 
                           N130);
   U2236 : AND2_X1 port map( A1 => regs_nxt_28_12_port, A2 => n27015, ZN => 
                           N131);
   U2237 : AND2_X1 port map( A1 => regs_nxt_28_13_port, A2 => n27015, ZN => 
                           N132);
   U2238 : AND2_X1 port map( A1 => regs_nxt_28_14_port, A2 => n27015, ZN => 
                           N133);
   U2239 : AND2_X1 port map( A1 => regs_nxt_28_15_port, A2 => n27016, ZN => 
                           N134);
   U2240 : AND2_X1 port map( A1 => regs_nxt_28_16_port, A2 => n27016, ZN => 
                           N135);
   U2241 : AND2_X1 port map( A1 => regs_nxt_28_17_port, A2 => n27016, ZN => 
                           N136);
   U2242 : AND2_X1 port map( A1 => regs_nxt_28_18_port, A2 => n27016, ZN => 
                           N137);
   U2243 : AND2_X1 port map( A1 => regs_nxt_28_19_port, A2 => n27016, ZN => 
                           N138);
   U2244 : AND2_X1 port map( A1 => regs_nxt_28_20_port, A2 => n27016, ZN => 
                           N139);
   U2245 : AND2_X1 port map( A1 => regs_nxt_28_21_port, A2 => n27016, ZN => 
                           N140);
   U2246 : AND2_X1 port map( A1 => regs_nxt_28_22_port, A2 => n27016, ZN => 
                           N141);
   U2247 : AND2_X1 port map( A1 => regs_nxt_28_23_port, A2 => n27016, ZN => 
                           N142);
   U2248 : AND2_X1 port map( A1 => regs_nxt_28_24_port, A2 => n27016, ZN => 
                           N143);
   U2249 : AND2_X1 port map( A1 => regs_nxt_28_25_port, A2 => n27016, ZN => 
                           N144);
   U2250 : AND2_X1 port map( A1 => regs_nxt_28_26_port, A2 => n27016, ZN => 
                           N145);
   U2251 : AND2_X1 port map( A1 => regs_nxt_28_27_port, A2 => n27016, ZN => 
                           N146);
   U2252 : AND2_X1 port map( A1 => regs_nxt_28_28_port, A2 => n27016, ZN => 
                           N147);
   U2253 : AND2_X1 port map( A1 => regs_nxt_28_29_port, A2 => n27016, ZN => 
                           N148);
   U2254 : AND2_X1 port map( A1 => regs_nxt_28_30_port, A2 => n27016, ZN => 
                           N149);
   U2255 : AND2_X1 port map( A1 => regs_nxt_28_31_port, A2 => n27016, ZN => 
                           N150);
   U2256 : AND2_X1 port map( A1 => regs_nxt_27_0_port, A2 => n27016, ZN => N151
                           );
   U2257 : AND2_X1 port map( A1 => regs_nxt_27_1_port, A2 => n27017, ZN => N152
                           );
   U2258 : AND2_X1 port map( A1 => regs_nxt_27_2_port, A2 => n27017, ZN => N153
                           );
   U2259 : AND2_X1 port map( A1 => regs_nxt_27_3_port, A2 => n27017, ZN => N154
                           );
   U2260 : AND2_X1 port map( A1 => regs_nxt_27_4_port, A2 => n27017, ZN => N155
                           );
   U2261 : AND2_X1 port map( A1 => regs_nxt_27_5_port, A2 => n27017, ZN => N156
                           );
   U2262 : AND2_X1 port map( A1 => regs_nxt_27_6_port, A2 => n27017, ZN => N157
                           );
   U2263 : AND2_X1 port map( A1 => regs_nxt_27_7_port, A2 => n27017, ZN => N158
                           );
   U2264 : AND2_X1 port map( A1 => regs_nxt_27_8_port, A2 => n27017, ZN => N159
                           );
   U2265 : AND2_X1 port map( A1 => regs_nxt_27_9_port, A2 => n27017, ZN => N160
                           );
   U2266 : AND2_X1 port map( A1 => regs_nxt_27_10_port, A2 => n27017, ZN => 
                           N161);
   U2267 : AND2_X1 port map( A1 => regs_nxt_27_11_port, A2 => n27017, ZN => 
                           N162);
   U2268 : AND2_X1 port map( A1 => regs_nxt_27_12_port, A2 => n27017, ZN => 
                           N163);
   U2269 : AND2_X1 port map( A1 => regs_nxt_27_13_port, A2 => n27017, ZN => 
                           N164);
   U2270 : AND2_X1 port map( A1 => regs_nxt_27_14_port, A2 => n27017, ZN => 
                           N165);
   U2271 : AND2_X1 port map( A1 => regs_nxt_27_15_port, A2 => n27017, ZN => 
                           N166);
   U2272 : AND2_X1 port map( A1 => regs_nxt_27_16_port, A2 => n27017, ZN => 
                           N167);
   U2273 : AND2_X1 port map( A1 => regs_nxt_27_17_port, A2 => n27017, ZN => 
                           N168);
   U2274 : AND2_X1 port map( A1 => regs_nxt_27_18_port, A2 => n27017, ZN => 
                           N169);
   U2275 : AND2_X1 port map( A1 => regs_nxt_27_19_port, A2 => n27018, ZN => 
                           N170);
   U2276 : AND2_X1 port map( A1 => regs_nxt_27_20_port, A2 => n27018, ZN => 
                           N171);
   U2277 : AND2_X1 port map( A1 => regs_nxt_27_21_port, A2 => n27018, ZN => 
                           N172);
   U2278 : AND2_X1 port map( A1 => regs_nxt_27_22_port, A2 => n27018, ZN => 
                           N173);
   U2279 : AND2_X1 port map( A1 => regs_nxt_27_23_port, A2 => n27018, ZN => 
                           N174);
   U2280 : AND2_X1 port map( A1 => regs_nxt_27_24_port, A2 => n27018, ZN => 
                           N175);
   U2281 : AND2_X1 port map( A1 => regs_nxt_27_25_port, A2 => n27018, ZN => 
                           N176);
   U2282 : AND2_X1 port map( A1 => regs_nxt_27_26_port, A2 => n27018, ZN => 
                           N177);
   U2283 : AND2_X1 port map( A1 => regs_nxt_27_27_port, A2 => n27018, ZN => 
                           N178);
   U2284 : AND2_X1 port map( A1 => regs_nxt_27_28_port, A2 => n27018, ZN => 
                           N179);
   U2285 : AND2_X1 port map( A1 => regs_nxt_27_29_port, A2 => n27018, ZN => 
                           N180);
   U2286 : AND2_X1 port map( A1 => regs_nxt_27_30_port, A2 => n27018, ZN => 
                           N181);
   U2287 : AND2_X1 port map( A1 => regs_nxt_27_31_port, A2 => n27018, ZN => 
                           N182);
   U2288 : AND2_X1 port map( A1 => regs_nxt_26_0_port, A2 => n27018, ZN => N183
                           );
   U2289 : AND2_X1 port map( A1 => regs_nxt_26_1_port, A2 => n27018, ZN => N184
                           );
   U2290 : AND2_X1 port map( A1 => regs_nxt_26_2_port, A2 => n27018, ZN => N185
                           );
   U2291 : AND2_X1 port map( A1 => regs_nxt_26_3_port, A2 => n27007, ZN => N186
                           );
   U2292 : AND2_X1 port map( A1 => regs_nxt_26_4_port, A2 => n27004, ZN => N187
                           );
   U2293 : AND2_X1 port map( A1 => regs_nxt_26_5_port, A2 => n27004, ZN => N188
                           );
   U2294 : AND2_X1 port map( A1 => regs_nxt_26_6_port, A2 => n27004, ZN => N189
                           );
   U2295 : AND2_X1 port map( A1 => regs_nxt_26_7_port, A2 => n27004, ZN => N190
                           );
   U2296 : AND2_X1 port map( A1 => regs_nxt_26_8_port, A2 => n27004, ZN => N191
                           );
   U2297 : AND2_X1 port map( A1 => regs_nxt_26_9_port, A2 => n27004, ZN => N192
                           );
   U2298 : AND2_X1 port map( A1 => regs_nxt_26_10_port, A2 => n27004, ZN => 
                           N193);
   U2299 : AND2_X1 port map( A1 => regs_nxt_26_11_port, A2 => n27004, ZN => 
                           N194);
   U2300 : AND2_X1 port map( A1 => regs_nxt_26_12_port, A2 => n27004, ZN => 
                           N195);
   U2301 : AND2_X1 port map( A1 => regs_nxt_26_13_port, A2 => n27004, ZN => 
                           N196);
   U2302 : AND2_X1 port map( A1 => regs_nxt_26_14_port, A2 => n27004, ZN => 
                           N197);
   U2303 : AND2_X1 port map( A1 => regs_nxt_26_15_port, A2 => n27004, ZN => 
                           N198);
   U2304 : AND2_X1 port map( A1 => regs_nxt_26_16_port, A2 => n27004, ZN => 
                           N199);
   U2305 : AND2_X1 port map( A1 => regs_nxt_26_17_port, A2 => n27005, ZN => 
                           N200);
   U2306 : AND2_X1 port map( A1 => regs_nxt_26_18_port, A2 => n27005, ZN => 
                           N201);
   U2307 : AND2_X1 port map( A1 => regs_nxt_26_19_port, A2 => n27005, ZN => 
                           N202);
   U2308 : AND2_X1 port map( A1 => regs_nxt_26_20_port, A2 => n27005, ZN => 
                           N203);
   U2309 : AND2_X1 port map( A1 => regs_nxt_26_21_port, A2 => n27005, ZN => 
                           N204);
   U2310 : AND2_X1 port map( A1 => regs_nxt_26_22_port, A2 => n27005, ZN => 
                           N205);
   U2311 : AND2_X1 port map( A1 => regs_nxt_26_23_port, A2 => n27005, ZN => 
                           N206);
   U2312 : AND2_X1 port map( A1 => regs_nxt_26_24_port, A2 => n27005, ZN => 
                           N207);
   U2313 : AND2_X1 port map( A1 => regs_nxt_26_25_port, A2 => n27005, ZN => 
                           N208);
   U2314 : AND2_X1 port map( A1 => regs_nxt_26_26_port, A2 => n27005, ZN => 
                           N209);
   U2315 : AND2_X1 port map( A1 => regs_nxt_26_27_port, A2 => n27005, ZN => 
                           N210);
   U2316 : AND2_X1 port map( A1 => regs_nxt_26_28_port, A2 => n27005, ZN => 
                           N211);
   U2317 : AND2_X1 port map( A1 => regs_nxt_26_29_port, A2 => n27005, ZN => 
                           N212);
   U2318 : AND2_X1 port map( A1 => regs_nxt_26_30_port, A2 => n27005, ZN => 
                           N213);
   U2319 : AND2_X1 port map( A1 => regs_nxt_26_31_port, A2 => n27005, ZN => 
                           N214);
   U2320 : AND2_X1 port map( A1 => regs_nxt_25_0_port, A2 => n27005, ZN => N215
                           );
   U2321 : AND2_X1 port map( A1 => regs_nxt_25_1_port, A2 => n27005, ZN => N216
                           );
   U2322 : AND2_X1 port map( A1 => regs_nxt_25_2_port, A2 => n27005, ZN => N217
                           );
   U2323 : AND2_X1 port map( A1 => regs_nxt_25_3_port, A2 => n27006, ZN => N218
                           );
   U2324 : AND2_X1 port map( A1 => regs_nxt_25_4_port, A2 => n27006, ZN => N219
                           );
   U2325 : AND2_X1 port map( A1 => regs_nxt_25_5_port, A2 => n27006, ZN => N220
                           );
   U2326 : AND2_X1 port map( A1 => regs_nxt_25_6_port, A2 => n27006, ZN => N221
                           );
   U2327 : AND2_X1 port map( A1 => regs_nxt_25_7_port, A2 => n27006, ZN => N222
                           );
   U2328 : AND2_X1 port map( A1 => regs_nxt_25_8_port, A2 => n27006, ZN => N223
                           );
   U2329 : AND2_X1 port map( A1 => regs_nxt_25_9_port, A2 => n27006, ZN => N224
                           );
   U2330 : AND2_X1 port map( A1 => regs_nxt_25_10_port, A2 => n27006, ZN => 
                           N225);
   U2331 : AND2_X1 port map( A1 => regs_nxt_25_11_port, A2 => n27006, ZN => 
                           N226);
   U2332 : AND2_X1 port map( A1 => regs_nxt_25_12_port, A2 => n27006, ZN => 
                           N227);
   U2333 : AND2_X1 port map( A1 => regs_nxt_25_13_port, A2 => n27006, ZN => 
                           N228);
   U2334 : AND2_X1 port map( A1 => regs_nxt_25_14_port, A2 => n27006, ZN => 
                           N229);
   U2335 : AND2_X1 port map( A1 => regs_nxt_25_15_port, A2 => n27006, ZN => 
                           N230);
   U2336 : AND2_X1 port map( A1 => regs_nxt_25_16_port, A2 => n27006, ZN => 
                           N231);
   U2337 : AND2_X1 port map( A1 => regs_nxt_25_17_port, A2 => n27006, ZN => 
                           N232);
   U2338 : AND2_X1 port map( A1 => regs_nxt_25_18_port, A2 => n27006, ZN => 
                           N233);
   U2339 : AND2_X1 port map( A1 => regs_nxt_25_19_port, A2 => n27006, ZN => 
                           N234);
   U2340 : AND2_X1 port map( A1 => regs_nxt_25_20_port, A2 => n27007, ZN => 
                           N235);
   U2341 : AND2_X1 port map( A1 => regs_nxt_25_21_port, A2 => n27007, ZN => 
                           N236);
   U2342 : AND2_X1 port map( A1 => regs_nxt_25_22_port, A2 => n27007, ZN => 
                           N237);
   U2343 : AND2_X1 port map( A1 => regs_nxt_25_23_port, A2 => n27007, ZN => 
                           N238);
   U2344 : AND2_X1 port map( A1 => regs_nxt_25_24_port, A2 => n27007, ZN => 
                           N239);
   U2345 : AND2_X1 port map( A1 => regs_nxt_25_25_port, A2 => n27007, ZN => 
                           N240);
   U2346 : AND2_X1 port map( A1 => regs_nxt_25_26_port, A2 => n27007, ZN => 
                           N241);
   U2347 : AND2_X1 port map( A1 => regs_nxt_25_27_port, A2 => n27007, ZN => 
                           N242);
   U2348 : AND2_X1 port map( A1 => regs_nxt_25_28_port, A2 => n27007, ZN => 
                           N243);
   U2349 : AND2_X1 port map( A1 => regs_nxt_25_29_port, A2 => n27007, ZN => 
                           N244);
   U2350 : AND2_X1 port map( A1 => regs_nxt_25_30_port, A2 => n27007, ZN => 
                           N245);
   U2351 : AND2_X1 port map( A1 => regs_nxt_25_31_port, A2 => n27007, ZN => 
                           N246);
   U2352 : AND2_X1 port map( A1 => regs_nxt_24_0_port, A2 => n27007, ZN => N247
                           );
   U2353 : AND2_X1 port map( A1 => regs_nxt_24_1_port, A2 => n27007, ZN => N248
                           );
   U2354 : AND2_X1 port map( A1 => regs_nxt_24_2_port, A2 => n27007, ZN => N249
                           );
   U2355 : AND2_X1 port map( A1 => regs_nxt_24_3_port, A2 => n27008, ZN => N250
                           );
   U2356 : AND2_X1 port map( A1 => regs_nxt_24_4_port, A2 => n27008, ZN => N251
                           );
   U2357 : AND2_X1 port map( A1 => regs_nxt_24_5_port, A2 => n27008, ZN => N252
                           );
   U2358 : AND2_X1 port map( A1 => regs_nxt_24_6_port, A2 => n27008, ZN => N253
                           );
   U2359 : AND2_X1 port map( A1 => regs_nxt_24_7_port, A2 => n27008, ZN => N254
                           );
   U2360 : AND2_X1 port map( A1 => regs_nxt_24_8_port, A2 => n27008, ZN => N255
                           );
   U2361 : AND2_X1 port map( A1 => regs_nxt_24_9_port, A2 => n27008, ZN => N256
                           );
   U2362 : AND2_X1 port map( A1 => regs_nxt_24_10_port, A2 => n27008, ZN => 
                           N257);
   U2363 : AND2_X1 port map( A1 => regs_nxt_24_11_port, A2 => n27008, ZN => 
                           N258);
   U2364 : AND2_X1 port map( A1 => regs_nxt_24_12_port, A2 => n27008, ZN => 
                           N259);
   U2365 : AND2_X1 port map( A1 => regs_nxt_24_13_port, A2 => n27008, ZN => 
                           N260);
   U2366 : AND2_X1 port map( A1 => regs_nxt_24_14_port, A2 => n27008, ZN => 
                           N261);
   U2367 : AND2_X1 port map( A1 => regs_nxt_24_15_port, A2 => n27008, ZN => 
                           N262);
   U2368 : AND2_X1 port map( A1 => regs_nxt_24_16_port, A2 => n27008, ZN => 
                           N263);
   U2369 : AND2_X1 port map( A1 => regs_nxt_24_17_port, A2 => n27008, ZN => 
                           N264);
   U2370 : AND2_X1 port map( A1 => regs_nxt_24_18_port, A2 => n27008, ZN => 
                           N265);
   U2371 : AND2_X1 port map( A1 => regs_nxt_24_19_port, A2 => n27008, ZN => 
                           N266);
   U2372 : AND2_X1 port map( A1 => regs_nxt_24_20_port, A2 => n27009, ZN => 
                           N267);
   U2373 : AND2_X1 port map( A1 => regs_nxt_24_21_port, A2 => n27009, ZN => 
                           N268);
   U2374 : AND2_X1 port map( A1 => regs_nxt_24_22_port, A2 => n27009, ZN => 
                           N269);
   U2375 : AND2_X1 port map( A1 => regs_nxt_24_23_port, A2 => n27009, ZN => 
                           N270);
   U2376 : AND2_X1 port map( A1 => regs_nxt_24_24_port, A2 => n27009, ZN => 
                           N271);
   U2377 : AND2_X1 port map( A1 => regs_nxt_24_25_port, A2 => n27009, ZN => 
                           N272);
   U2378 : AND2_X1 port map( A1 => regs_nxt_24_26_port, A2 => n27009, ZN => 
                           N273);
   U2379 : AND2_X1 port map( A1 => regs_nxt_24_27_port, A2 => n27009, ZN => 
                           N274);
   U2380 : AND2_X1 port map( A1 => regs_nxt_24_28_port, A2 => n27009, ZN => 
                           N275);
   U2381 : AND2_X1 port map( A1 => regs_nxt_24_29_port, A2 => n27009, ZN => 
                           N276);
   U2382 : AND2_X1 port map( A1 => regs_nxt_24_30_port, A2 => n27009, ZN => 
                           N277);
   U2383 : AND2_X1 port map( A1 => regs_nxt_24_31_port, A2 => n27009, ZN => 
                           N278);
   U2384 : AND2_X1 port map( A1 => regs_nxt_23_0_port, A2 => n27009, ZN => N279
                           );
   U2385 : AND2_X1 port map( A1 => regs_nxt_23_1_port, A2 => n27009, ZN => N280
                           );
   U2386 : AND2_X1 port map( A1 => regs_nxt_23_2_port, A2 => n27009, ZN => N281
                           );
   U2387 : AND2_X1 port map( A1 => regs_nxt_23_3_port, A2 => n27009, ZN => N282
                           );
   U2388 : AND2_X1 port map( A1 => regs_nxt_23_4_port, A2 => n27010, ZN => N283
                           );
   U2389 : AND2_X1 port map( A1 => regs_nxt_23_5_port, A2 => n27010, ZN => N284
                           );
   U2390 : AND2_X1 port map( A1 => regs_nxt_23_6_port, A2 => n27010, ZN => N285
                           );
   U2391 : AND2_X1 port map( A1 => regs_nxt_23_7_port, A2 => n27010, ZN => N286
                           );
   U2392 : AND2_X1 port map( A1 => regs_nxt_23_8_port, A2 => n27010, ZN => N287
                           );
   U2393 : AND2_X1 port map( A1 => regs_nxt_23_9_port, A2 => n27010, ZN => N288
                           );
   U2394 : AND2_X1 port map( A1 => regs_nxt_23_10_port, A2 => n27010, ZN => 
                           N289);
   U2395 : AND2_X1 port map( A1 => regs_nxt_23_11_port, A2 => n27010, ZN => 
                           N290);
   U2396 : AND2_X1 port map( A1 => regs_nxt_23_12_port, A2 => n27010, ZN => 
                           N291);
   U2397 : AND2_X1 port map( A1 => regs_nxt_23_13_port, A2 => n27010, ZN => 
                           N292);
   U2398 : AND2_X1 port map( A1 => regs_nxt_23_14_port, A2 => n27010, ZN => 
                           N293);
   U2399 : AND2_X1 port map( A1 => regs_nxt_23_15_port, A2 => n27010, ZN => 
                           N294);
   U2400 : AND2_X1 port map( A1 => regs_nxt_23_16_port, A2 => n27010, ZN => 
                           N295);
   U2401 : AND2_X1 port map( A1 => regs_nxt_23_17_port, A2 => n27010, ZN => 
                           N296);
   U2402 : AND2_X1 port map( A1 => regs_nxt_23_18_port, A2 => n27010, ZN => 
                           N297);
   U2403 : AND2_X1 port map( A1 => regs_nxt_23_19_port, A2 => n27010, ZN => 
                           N298);
   U2404 : AND2_X1 port map( A1 => regs_nxt_23_20_port, A2 => n27010, ZN => 
                           N299);
   U2405 : AND2_X1 port map( A1 => regs_nxt_23_21_port, A2 => n27011, ZN => 
                           N300);
   U2406 : AND2_X1 port map( A1 => regs_nxt_23_22_port, A2 => n27011, ZN => 
                           N301);
   U2407 : AND2_X1 port map( A1 => regs_nxt_23_23_port, A2 => n27011, ZN => 
                           N302);
   U2408 : AND2_X1 port map( A1 => regs_nxt_23_24_port, A2 => n27011, ZN => 
                           N303);
   U2409 : AND2_X1 port map( A1 => regs_nxt_23_25_port, A2 => n27011, ZN => 
                           N304);
   U2410 : AND2_X1 port map( A1 => regs_nxt_23_26_port, A2 => n27011, ZN => 
                           N305);
   U2411 : AND2_X1 port map( A1 => regs_nxt_23_27_port, A2 => n27011, ZN => 
                           N306);
   U2412 : AND2_X1 port map( A1 => regs_nxt_23_28_port, A2 => n27011, ZN => 
                           N307);
   U2413 : AND2_X1 port map( A1 => regs_nxt_23_29_port, A2 => n27011, ZN => 
                           N308);
   U2414 : AND2_X1 port map( A1 => regs_nxt_23_30_port, A2 => n27011, ZN => 
                           N309);
   U2415 : AND2_X1 port map( A1 => regs_nxt_23_31_port, A2 => n27026, ZN => 
                           N310);
   U2416 : AND2_X1 port map( A1 => regs_nxt_22_0_port, A2 => n27026, ZN => N311
                           );
   U2417 : AND2_X1 port map( A1 => regs_nxt_22_1_port, A2 => n27026, ZN => N312
                           );
   U2418 : AND2_X1 port map( A1 => regs_nxt_22_2_port, A2 => n27026, ZN => N313
                           );
   U2419 : AND2_X1 port map( A1 => regs_nxt_22_3_port, A2 => n27026, ZN => N314
                           );
   U2420 : AND2_X1 port map( A1 => regs_nxt_22_4_port, A2 => n27026, ZN => N315
                           );
   U2421 : AND2_X1 port map( A1 => regs_nxt_22_5_port, A2 => n27026, ZN => N316
                           );
   U2422 : AND2_X1 port map( A1 => regs_nxt_22_6_port, A2 => n27026, ZN => N317
                           );
   U2423 : AND2_X1 port map( A1 => regs_nxt_22_7_port, A2 => n27026, ZN => N318
                           );
   U2424 : AND2_X1 port map( A1 => regs_nxt_22_8_port, A2 => n27026, ZN => N319
                           );
   U2425 : AND2_X1 port map( A1 => regs_nxt_22_9_port, A2 => n27026, ZN => N320
                           );
   U2426 : AND2_X1 port map( A1 => regs_nxt_22_10_port, A2 => n27026, ZN => 
                           N321);
   U2427 : AND2_X1 port map( A1 => regs_nxt_22_11_port, A2 => n27027, ZN => 
                           N322);
   U2428 : AND2_X1 port map( A1 => regs_nxt_22_12_port, A2 => n27027, ZN => 
                           N323);
   U2429 : AND2_X1 port map( A1 => regs_nxt_22_13_port, A2 => n27027, ZN => 
                           N324);
   U2430 : AND2_X1 port map( A1 => regs_nxt_22_14_port, A2 => n27027, ZN => 
                           N325);
   U2431 : AND2_X1 port map( A1 => regs_nxt_22_15_port, A2 => n27027, ZN => 
                           N326);
   U2432 : AND2_X1 port map( A1 => regs_nxt_22_16_port, A2 => n27027, ZN => 
                           N327);
   U2433 : AND2_X1 port map( A1 => regs_nxt_22_17_port, A2 => n27027, ZN => 
                           N328);
   U2434 : AND2_X1 port map( A1 => regs_nxt_22_18_port, A2 => n27027, ZN => 
                           N329);
   U2435 : AND2_X1 port map( A1 => regs_nxt_22_19_port, A2 => n27027, ZN => 
                           N330);
   U2436 : AND2_X1 port map( A1 => regs_nxt_22_20_port, A2 => n27027, ZN => 
                           N331);
   U2437 : AND2_X1 port map( A1 => regs_nxt_22_21_port, A2 => n27027, ZN => 
                           N332);
   U2438 : AND2_X1 port map( A1 => regs_nxt_22_22_port, A2 => n27027, ZN => 
                           N333);
   U2439 : AND2_X1 port map( A1 => regs_nxt_22_23_port, A2 => n27027, ZN => 
                           N334);
   U2440 : AND2_X1 port map( A1 => regs_nxt_22_24_port, A2 => n27027, ZN => 
                           N335);
   U2441 : AND2_X1 port map( A1 => regs_nxt_22_25_port, A2 => n27027, ZN => 
                           N336);
   U2442 : AND2_X1 port map( A1 => regs_nxt_22_26_port, A2 => n27027, ZN => 
                           N337);
   U2443 : AND2_X1 port map( A1 => regs_nxt_22_27_port, A2 => n27027, ZN => 
                           N338);
   U2444 : AND2_X1 port map( A1 => regs_nxt_22_28_port, A2 => n27028, ZN => 
                           N339);
   U2445 : AND2_X1 port map( A1 => regs_nxt_22_29_port, A2 => n27028, ZN => 
                           N340);
   U2446 : AND2_X1 port map( A1 => regs_nxt_22_30_port, A2 => n27028, ZN => 
                           N341);
   U2447 : AND2_X1 port map( A1 => regs_nxt_22_31_port, A2 => n27028, ZN => 
                           N342);
   U2448 : AND2_X1 port map( A1 => regs_nxt_21_0_port, A2 => n27028, ZN => N343
                           );
   U2449 : AND2_X1 port map( A1 => regs_nxt_21_1_port, A2 => n27028, ZN => N344
                           );
   U2450 : AND2_X1 port map( A1 => regs_nxt_21_2_port, A2 => n27028, ZN => N345
                           );
   U2451 : AND2_X1 port map( A1 => regs_nxt_21_3_port, A2 => n27028, ZN => N346
                           );
   U2452 : AND2_X1 port map( A1 => regs_nxt_21_4_port, A2 => n27028, ZN => N347
                           );
   U2453 : AND2_X1 port map( A1 => regs_nxt_21_5_port, A2 => n27028, ZN => N348
                           );
   U2454 : AND2_X1 port map( A1 => regs_nxt_21_6_port, A2 => n27028, ZN => N349
                           );
   U2455 : AND2_X1 port map( A1 => regs_nxt_21_7_port, A2 => n27028, ZN => N350
                           );
   U2456 : AND2_X1 port map( A1 => regs_nxt_21_8_port, A2 => n27028, ZN => N351
                           );
   U2457 : AND2_X1 port map( A1 => regs_nxt_21_9_port, A2 => n27028, ZN => N352
                           );
   U2458 : AND2_X1 port map( A1 => regs_nxt_21_10_port, A2 => n27028, ZN => 
                           N353);
   U2459 : AND2_X1 port map( A1 => regs_nxt_21_11_port, A2 => n27028, ZN => 
                           N354);
   U2460 : AND2_X1 port map( A1 => regs_nxt_21_12_port, A2 => n27029, ZN => 
                           N355);
   U2461 : AND2_X1 port map( A1 => regs_nxt_21_13_port, A2 => n27029, ZN => 
                           N356);
   U2462 : AND2_X1 port map( A1 => regs_nxt_21_14_port, A2 => n27029, ZN => 
                           N357);
   U2463 : AND2_X1 port map( A1 => regs_nxt_21_15_port, A2 => n27029, ZN => 
                           N358);
   U2464 : AND2_X1 port map( A1 => regs_nxt_21_16_port, A2 => n27029, ZN => 
                           N359);
   U2465 : AND2_X1 port map( A1 => regs_nxt_21_17_port, A2 => n27029, ZN => 
                           N360);
   U2466 : AND2_X1 port map( A1 => regs_nxt_21_18_port, A2 => n27029, ZN => 
                           N361);
   U2467 : AND2_X1 port map( A1 => regs_nxt_21_19_port, A2 => n27029, ZN => 
                           N362);
   U2468 : AND2_X1 port map( A1 => regs_nxt_21_20_port, A2 => n27029, ZN => 
                           N363);
   U2469 : AND2_X1 port map( A1 => regs_nxt_21_21_port, A2 => n27029, ZN => 
                           N364);
   U2470 : AND2_X1 port map( A1 => regs_nxt_21_22_port, A2 => n27029, ZN => 
                           N365);
   U2471 : AND2_X1 port map( A1 => regs_nxt_21_23_port, A2 => n27029, ZN => 
                           N366);
   U2472 : AND2_X1 port map( A1 => regs_nxt_21_24_port, A2 => n27029, ZN => 
                           N367);
   U2473 : AND2_X1 port map( A1 => regs_nxt_21_25_port, A2 => n27029, ZN => 
                           N368);
   U2474 : AND2_X1 port map( A1 => regs_nxt_21_26_port, A2 => n27029, ZN => 
                           N369);
   U2475 : AND2_X1 port map( A1 => regs_nxt_21_27_port, A2 => n27030, ZN => 
                           N370);
   U2476 : AND2_X1 port map( A1 => regs_nxt_21_28_port, A2 => n27030, ZN => 
                           N371);
   U2477 : AND2_X1 port map( A1 => regs_nxt_21_29_port, A2 => n27030, ZN => 
                           N372);
   U2478 : AND2_X1 port map( A1 => regs_nxt_21_30_port, A2 => n27030, ZN => 
                           N373);
   U2479 : AND2_X1 port map( A1 => regs_nxt_21_31_port, A2 => n27030, ZN => 
                           N374);
   U2480 : AND2_X1 port map( A1 => regs_nxt_20_0_port, A2 => n27030, ZN => N375
                           );
   U2481 : AND2_X1 port map( A1 => regs_nxt_20_1_port, A2 => n27030, ZN => N376
                           );
   U2482 : AND2_X1 port map( A1 => regs_nxt_20_2_port, A2 => n27030, ZN => N377
                           );
   U2483 : AND2_X1 port map( A1 => regs_nxt_20_3_port, A2 => n27030, ZN => N378
                           );
   U2484 : AND2_X1 port map( A1 => regs_nxt_20_4_port, A2 => n27030, ZN => N379
                           );
   U2485 : AND2_X1 port map( A1 => regs_nxt_20_5_port, A2 => n27030, ZN => N380
                           );
   U2486 : AND2_X1 port map( A1 => regs_nxt_20_6_port, A2 => n27030, ZN => N381
                           );
   U2487 : AND2_X1 port map( A1 => regs_nxt_20_7_port, A2 => n27030, ZN => N382
                           );
   U2488 : AND2_X1 port map( A1 => regs_nxt_20_8_port, A2 => n27030, ZN => N383
                           );
   U2489 : AND2_X1 port map( A1 => regs_nxt_20_9_port, A2 => n27030, ZN => N384
                           );
   U2490 : AND2_X1 port map( A1 => regs_nxt_20_10_port, A2 => n27030, ZN => 
                           N385);
   U2491 : AND2_X1 port map( A1 => regs_nxt_20_11_port, A2 => n27030, ZN => 
                           N386);
   U2492 : AND2_X1 port map( A1 => regs_nxt_20_12_port, A2 => n27031, ZN => 
                           N387);
   U2493 : AND2_X1 port map( A1 => regs_nxt_20_13_port, A2 => n27031, ZN => 
                           N388);
   U2494 : AND2_X1 port map( A1 => regs_nxt_20_14_port, A2 => n27031, ZN => 
                           N389);
   U2495 : AND2_X1 port map( A1 => regs_nxt_20_15_port, A2 => n27031, ZN => 
                           N390);
   U2496 : AND2_X1 port map( A1 => regs_nxt_20_16_port, A2 => n27031, ZN => 
                           N391);
   U2497 : AND2_X1 port map( A1 => regs_nxt_20_17_port, A2 => n27031, ZN => 
                           N392);
   U2498 : AND2_X1 port map( A1 => regs_nxt_20_18_port, A2 => n27031, ZN => 
                           N393);
   U2499 : AND2_X1 port map( A1 => regs_nxt_20_19_port, A2 => n27031, ZN => 
                           N394);
   U2500 : AND2_X1 port map( A1 => regs_nxt_20_20_port, A2 => n27031, ZN => 
                           N395);
   U2501 : AND2_X1 port map( A1 => regs_nxt_20_21_port, A2 => n27031, ZN => 
                           N396);
   U2502 : AND2_X1 port map( A1 => regs_nxt_20_22_port, A2 => n27031, ZN => 
                           N397);
   U2503 : AND2_X1 port map( A1 => regs_nxt_20_23_port, A2 => n27031, ZN => 
                           N398);
   U2504 : AND2_X1 port map( A1 => regs_nxt_20_24_port, A2 => n27031, ZN => 
                           N399);
   U2505 : AND2_X1 port map( A1 => regs_nxt_20_25_port, A2 => n27031, ZN => 
                           N400);
   U2506 : AND2_X1 port map( A1 => regs_nxt_20_26_port, A2 => n27031, ZN => 
                           N401);
   U2507 : AND2_X1 port map( A1 => regs_nxt_20_27_port, A2 => n27031, ZN => 
                           N402);
   U2508 : AND2_X1 port map( A1 => regs_nxt_20_28_port, A2 => n27032, ZN => 
                           N403);
   U2509 : AND2_X1 port map( A1 => regs_nxt_20_29_port, A2 => n27032, ZN => 
                           N404);
   U2510 : AND2_X1 port map( A1 => regs_nxt_20_30_port, A2 => n27032, ZN => 
                           N405);
   U2511 : AND2_X1 port map( A1 => regs_nxt_20_31_port, A2 => n27032, ZN => 
                           N406);
   U2512 : AND2_X1 port map( A1 => regs_nxt_19_0_port, A2 => n27032, ZN => N407
                           );
   U2513 : AND2_X1 port map( A1 => regs_nxt_19_1_port, A2 => n27032, ZN => N408
                           );
   U2514 : AND2_X1 port map( A1 => regs_nxt_19_2_port, A2 => n27032, ZN => N409
                           );
   U2515 : AND2_X1 port map( A1 => regs_nxt_19_3_port, A2 => n27032, ZN => N410
                           );
   U2516 : AND2_X1 port map( A1 => regs_nxt_19_4_port, A2 => n27032, ZN => N411
                           );
   U2517 : AND2_X1 port map( A1 => regs_nxt_19_5_port, A2 => n27032, ZN => N412
                           );
   U2518 : AND2_X1 port map( A1 => regs_nxt_19_6_port, A2 => n27032, ZN => N413
                           );
   U2519 : AND2_X1 port map( A1 => regs_nxt_19_7_port, A2 => n27032, ZN => N414
                           );
   U2520 : AND2_X1 port map( A1 => regs_nxt_19_8_port, A2 => n27032, ZN => N415
                           );
   U2521 : AND2_X1 port map( A1 => regs_nxt_19_9_port, A2 => n27032, ZN => N416
                           );
   U2522 : AND2_X1 port map( A1 => regs_nxt_19_10_port, A2 => n27032, ZN => 
                           N417);
   U2523 : AND2_X1 port map( A1 => regs_nxt_19_11_port, A2 => n27032, ZN => 
                           N418);
   U2524 : AND2_X1 port map( A1 => regs_nxt_19_12_port, A2 => n27032, ZN => 
                           N419);
   U2525 : AND2_X1 port map( A1 => regs_nxt_19_13_port, A2 => n27033, ZN => 
                           N420);
   U2526 : AND2_X1 port map( A1 => regs_nxt_19_14_port, A2 => n27033, ZN => 
                           N421);
   U2527 : AND2_X1 port map( A1 => regs_nxt_19_15_port, A2 => n27033, ZN => 
                           N422);
   U2528 : AND2_X1 port map( A1 => regs_nxt_19_16_port, A2 => n27033, ZN => 
                           N423);
   U2529 : AND2_X1 port map( A1 => regs_nxt_19_17_port, A2 => n27033, ZN => 
                           N424);
   U2530 : AND2_X1 port map( A1 => regs_nxt_19_18_port, A2 => n27033, ZN => 
                           N425);
   U2531 : AND2_X1 port map( A1 => regs_nxt_19_19_port, A2 => n27033, ZN => 
                           N426);
   U2532 : AND2_X1 port map( A1 => regs_nxt_19_20_port, A2 => n27033, ZN => 
                           N427);
   U2533 : AND2_X1 port map( A1 => regs_nxt_19_21_port, A2 => n27033, ZN => 
                           N428);
   U2534 : AND2_X1 port map( A1 => regs_nxt_19_22_port, A2 => n27022, ZN => 
                           N429);
   U2535 : AND2_X1 port map( A1 => regs_nxt_19_23_port, A2 => n27019, ZN => 
                           N430);
   U2536 : AND2_X1 port map( A1 => regs_nxt_19_24_port, A2 => n27019, ZN => 
                           N431);
   U2537 : AND2_X1 port map( A1 => regs_nxt_19_25_port, A2 => n27019, ZN => 
                           N432);
   U2538 : AND2_X1 port map( A1 => regs_nxt_19_26_port, A2 => n27019, ZN => 
                           N433);
   U2539 : AND2_X1 port map( A1 => regs_nxt_19_27_port, A2 => n27019, ZN => 
                           N434);
   U2540 : AND2_X1 port map( A1 => regs_nxt_19_28_port, A2 => n27019, ZN => 
                           N435);
   U2541 : AND2_X1 port map( A1 => regs_nxt_19_29_port, A2 => n27019, ZN => 
                           N436);
   U2542 : AND2_X1 port map( A1 => regs_nxt_19_30_port, A2 => n27019, ZN => 
                           N437);
   U2543 : AND2_X1 port map( A1 => regs_nxt_19_31_port, A2 => n27019, ZN => 
                           N438);
   U2544 : AND2_X1 port map( A1 => regs_nxt_18_0_port, A2 => n27019, ZN => N439
                           );
   U2545 : AND2_X1 port map( A1 => regs_nxt_18_1_port, A2 => n27019, ZN => N440
                           );
   U2546 : AND2_X1 port map( A1 => regs_nxt_18_2_port, A2 => n27019, ZN => N441
                           );
   U2547 : AND2_X1 port map( A1 => regs_nxt_18_3_port, A2 => n27019, ZN => N442
                           );
   U2548 : AND2_X1 port map( A1 => regs_nxt_18_4_port, A2 => n27019, ZN => N443
                           );
   U2549 : AND2_X1 port map( A1 => regs_nxt_18_5_port, A2 => n27019, ZN => N444
                           );
   U2550 : AND2_X1 port map( A1 => regs_nxt_18_6_port, A2 => n27019, ZN => N445
                           );
   U2551 : AND2_X1 port map( A1 => regs_nxt_18_7_port, A2 => n27019, ZN => N446
                           );
   U2552 : AND2_X1 port map( A1 => regs_nxt_18_8_port, A2 => n27020, ZN => N447
                           );
   U2553 : AND2_X1 port map( A1 => regs_nxt_18_9_port, A2 => n27020, ZN => N448
                           );
   U2554 : AND2_X1 port map( A1 => regs_nxt_18_10_port, A2 => n27020, ZN => 
                           N449);
   U2555 : AND2_X1 port map( A1 => regs_nxt_18_11_port, A2 => n27020, ZN => 
                           N450);
   U2556 : AND2_X1 port map( A1 => regs_nxt_18_12_port, A2 => n27020, ZN => 
                           N451);
   U2557 : AND2_X1 port map( A1 => regs_nxt_18_13_port, A2 => n27020, ZN => 
                           N452);
   U2558 : AND2_X1 port map( A1 => regs_nxt_18_14_port, A2 => n27020, ZN => 
                           N453);
   U2559 : AND2_X1 port map( A1 => regs_nxt_18_15_port, A2 => n27020, ZN => 
                           N454);
   U2560 : AND2_X1 port map( A1 => regs_nxt_18_16_port, A2 => n27020, ZN => 
                           N455);
   U2561 : AND2_X1 port map( A1 => regs_nxt_18_17_port, A2 => n27020, ZN => 
                           N456);
   U2562 : AND2_X1 port map( A1 => regs_nxt_18_18_port, A2 => n27020, ZN => 
                           N457);
   U2563 : AND2_X1 port map( A1 => regs_nxt_18_19_port, A2 => n27020, ZN => 
                           N458);
   U2564 : AND2_X1 port map( A1 => regs_nxt_18_20_port, A2 => n27020, ZN => 
                           N459);
   U2565 : AND2_X1 port map( A1 => regs_nxt_18_21_port, A2 => n27020, ZN => 
                           N460);
   U2566 : AND2_X1 port map( A1 => regs_nxt_18_22_port, A2 => n27020, ZN => 
                           N461);
   U2567 : AND2_X1 port map( A1 => regs_nxt_18_23_port, A2 => n27020, ZN => 
                           N462);
   U2568 : AND2_X1 port map( A1 => regs_nxt_18_24_port, A2 => n27021, ZN => 
                           N463);
   U2569 : AND2_X1 port map( A1 => regs_nxt_18_25_port, A2 => n27021, ZN => 
                           N464);
   U2570 : AND2_X1 port map( A1 => regs_nxt_18_26_port, A2 => n27021, ZN => 
                           N465);
   U2571 : AND2_X1 port map( A1 => regs_nxt_18_27_port, A2 => n27021, ZN => 
                           N466);
   U2572 : AND2_X1 port map( A1 => regs_nxt_18_28_port, A2 => n27021, ZN => 
                           N467);
   U2573 : AND2_X1 port map( A1 => regs_nxt_18_29_port, A2 => n27021, ZN => 
                           N468);
   U2574 : AND2_X1 port map( A1 => regs_nxt_18_30_port, A2 => n27021, ZN => 
                           N469);
   U2575 : AND2_X1 port map( A1 => regs_nxt_18_31_port, A2 => n27021, ZN => 
                           N470);
   U2576 : AND2_X1 port map( A1 => regs_nxt_17_0_port, A2 => n27021, ZN => N471
                           );
   U2577 : AND2_X1 port map( A1 => regs_nxt_17_1_port, A2 => n27021, ZN => N472
                           );
   U2578 : AND2_X1 port map( A1 => regs_nxt_17_2_port, A2 => n27021, ZN => N473
                           );
   U2579 : AND2_X1 port map( A1 => regs_nxt_17_3_port, A2 => n27021, ZN => N474
                           );
   U2580 : AND2_X1 port map( A1 => regs_nxt_17_4_port, A2 => n27021, ZN => N475
                           );
   U2581 : AND2_X1 port map( A1 => regs_nxt_17_5_port, A2 => n27021, ZN => N476
                           );
   U2582 : AND2_X1 port map( A1 => regs_nxt_17_6_port, A2 => n27021, ZN => N477
                           );
   U2583 : AND2_X1 port map( A1 => regs_nxt_17_7_port, A2 => n27021, ZN => N478
                           );
   U2584 : AND2_X1 port map( A1 => regs_nxt_17_8_port, A2 => n27021, ZN => N479
                           );
   U2585 : AND2_X1 port map( A1 => regs_nxt_17_9_port, A2 => n27022, ZN => N480
                           );
   U2586 : AND2_X1 port map( A1 => regs_nxt_17_10_port, A2 => n27022, ZN => 
                           N481);
   U2587 : AND2_X1 port map( A1 => regs_nxt_17_11_port, A2 => n27022, ZN => 
                           N482);
   U2588 : AND2_X1 port map( A1 => regs_nxt_17_12_port, A2 => n27022, ZN => 
                           N483);
   U2589 : AND2_X1 port map( A1 => regs_nxt_17_13_port, A2 => n27022, ZN => 
                           N484);
   U2590 : AND2_X1 port map( A1 => regs_nxt_17_14_port, A2 => n27022, ZN => 
                           N485);
   U2591 : AND2_X1 port map( A1 => regs_nxt_17_15_port, A2 => n27022, ZN => 
                           N486);
   U2592 : AND2_X1 port map( A1 => regs_nxt_17_16_port, A2 => n27022, ZN => 
                           N487);
   U2593 : AND2_X1 port map( A1 => regs_nxt_17_17_port, A2 => n27022, ZN => 
                           N488);
   U2594 : AND2_X1 port map( A1 => regs_nxt_17_18_port, A2 => n27022, ZN => 
                           N489);
   U2595 : AND2_X1 port map( A1 => regs_nxt_17_19_port, A2 => n27022, ZN => 
                           N490);
   U2596 : AND2_X1 port map( A1 => regs_nxt_17_20_port, A2 => n27022, ZN => 
                           N491);
   U2597 : AND2_X1 port map( A1 => regs_nxt_17_21_port, A2 => n27022, ZN => 
                           N492);
   U2598 : AND2_X1 port map( A1 => regs_nxt_17_22_port, A2 => n27022, ZN => 
                           N493);
   U2599 : AND2_X1 port map( A1 => regs_nxt_17_23_port, A2 => n27022, ZN => 
                           N494);
   U2600 : AND2_X1 port map( A1 => regs_nxt_17_24_port, A2 => n27023, ZN => 
                           N495);
   U2601 : AND2_X1 port map( A1 => regs_nxt_17_25_port, A2 => n27023, ZN => 
                           N496);
   U2602 : AND2_X1 port map( A1 => regs_nxt_17_26_port, A2 => n27023, ZN => 
                           N497);
   U2603 : AND2_X1 port map( A1 => regs_nxt_17_27_port, A2 => n27023, ZN => 
                           N498);
   U2604 : AND2_X1 port map( A1 => regs_nxt_17_28_port, A2 => n27023, ZN => 
                           N499);
   U2605 : AND2_X1 port map( A1 => regs_nxt_17_29_port, A2 => n27023, ZN => 
                           N500);
   U2606 : AND2_X1 port map( A1 => regs_nxt_17_30_port, A2 => n27023, ZN => 
                           N501);
   U2607 : AND2_X1 port map( A1 => regs_nxt_17_31_port, A2 => n27023, ZN => 
                           N502);
   U2608 : AND2_X1 port map( A1 => regs_nxt_16_0_port, A2 => n27023, ZN => N503
                           );
   U2609 : AND2_X1 port map( A1 => regs_nxt_16_1_port, A2 => n27023, ZN => N504
                           );
   U2610 : AND2_X1 port map( A1 => regs_nxt_16_2_port, A2 => n27023, ZN => N505
                           );
   U2611 : AND2_X1 port map( A1 => regs_nxt_16_3_port, A2 => n27023, ZN => N506
                           );
   U2612 : AND2_X1 port map( A1 => regs_nxt_16_4_port, A2 => n27023, ZN => N507
                           );
   U2613 : AND2_X1 port map( A1 => regs_nxt_16_5_port, A2 => n27023, ZN => N508
                           );
   U2614 : AND2_X1 port map( A1 => regs_nxt_16_6_port, A2 => n27023, ZN => N509
                           );
   U2615 : AND2_X1 port map( A1 => regs_nxt_16_7_port, A2 => n27023, ZN => N510
                           );
   U2616 : AND2_X1 port map( A1 => regs_nxt_16_8_port, A2 => n27024, ZN => N511
                           );
   U2617 : AND2_X1 port map( A1 => regs_nxt_16_9_port, A2 => n27024, ZN => N512
                           );
   U2618 : AND2_X1 port map( A1 => regs_nxt_16_10_port, A2 => n27024, ZN => 
                           N513);
   U2619 : AND2_X1 port map( A1 => regs_nxt_16_11_port, A2 => n27024, ZN => 
                           N514);
   U2620 : AND2_X1 port map( A1 => regs_nxt_16_12_port, A2 => n27024, ZN => 
                           N515);
   U2621 : AND2_X1 port map( A1 => regs_nxt_16_13_port, A2 => n27024, ZN => 
                           N516);
   U2622 : AND2_X1 port map( A1 => regs_nxt_16_14_port, A2 => n27024, ZN => 
                           N517);
   U2623 : AND2_X1 port map( A1 => regs_nxt_16_15_port, A2 => n27024, ZN => 
                           N518);
   U2624 : AND2_X1 port map( A1 => regs_nxt_16_16_port, A2 => n27024, ZN => 
                           N519);
   U2625 : AND2_X1 port map( A1 => regs_nxt_16_17_port, A2 => n27024, ZN => 
                           N520);
   U2626 : AND2_X1 port map( A1 => regs_nxt_16_18_port, A2 => n27024, ZN => 
                           N521);
   U2627 : AND2_X1 port map( A1 => regs_nxt_16_19_port, A2 => n27024, ZN => 
                           N522);
   U2628 : AND2_X1 port map( A1 => regs_nxt_16_20_port, A2 => n27024, ZN => 
                           N523);
   U2629 : AND2_X1 port map( A1 => regs_nxt_16_21_port, A2 => n27024, ZN => 
                           N524);
   U2630 : AND2_X1 port map( A1 => regs_nxt_16_22_port, A2 => n27024, ZN => 
                           N525);
   U2631 : AND2_X1 port map( A1 => regs_nxt_16_23_port, A2 => n27024, ZN => 
                           N526);
   U2632 : AND2_X1 port map( A1 => regs_nxt_16_24_port, A2 => n27024, ZN => 
                           N527);
   U2633 : AND2_X1 port map( A1 => regs_nxt_16_25_port, A2 => n27025, ZN => 
                           N528);
   U2634 : AND2_X1 port map( A1 => regs_nxt_16_26_port, A2 => n27025, ZN => 
                           N529);
   U2635 : AND2_X1 port map( A1 => regs_nxt_16_27_port, A2 => n27025, ZN => 
                           N530);
   U2636 : AND2_X1 port map( A1 => regs_nxt_16_28_port, A2 => n27025, ZN => 
                           N531);
   U2637 : AND2_X1 port map( A1 => regs_nxt_16_29_port, A2 => n27025, ZN => 
                           N532);
   U2638 : AND2_X1 port map( A1 => regs_nxt_16_30_port, A2 => n27025, ZN => 
                           N533);
   U2639 : AND2_X1 port map( A1 => regs_nxt_16_31_port, A2 => n27025, ZN => 
                           N534);
   U2640 : AND2_X1 port map( A1 => regs_nxt_15_0_port, A2 => n27025, ZN => N535
                           );
   U2641 : AND2_X1 port map( A1 => regs_nxt_15_1_port, A2 => n27025, ZN => N536
                           );
   U2642 : AND2_X1 port map( A1 => regs_nxt_15_2_port, A2 => n27025, ZN => N537
                           );
   U2643 : AND2_X1 port map( A1 => regs_nxt_15_3_port, A2 => n27025, ZN => N538
                           );
   U2644 : AND2_X1 port map( A1 => regs_nxt_15_4_port, A2 => n27025, ZN => N539
                           );
   U2645 : AND2_X1 port map( A1 => regs_nxt_15_5_port, A2 => n27025, ZN => N540
                           );
   U2646 : AND2_X1 port map( A1 => regs_nxt_15_6_port, A2 => n27025, ZN => N541
                           );
   U2647 : AND2_X1 port map( A1 => regs_nxt_15_7_port, A2 => n27025, ZN => N542
                           );
   U2648 : AND2_X1 port map( A1 => regs_nxt_15_8_port, A2 => n27025, ZN => N543
                           );
   U2649 : AND2_X1 port map( A1 => regs_nxt_15_9_port, A2 => n27026, ZN => N544
                           );
   U2650 : AND2_X1 port map( A1 => regs_nxt_15_10_port, A2 => n27026, ZN => 
                           N545);
   U2651 : AND2_X1 port map( A1 => regs_nxt_15_11_port, A2 => n27026, ZN => 
                           N546);
   U2652 : AND2_X1 port map( A1 => regs_nxt_15_12_port, A2 => n27026, ZN => 
                           N547);
   U2653 : AND2_X1 port map( A1 => regs_nxt_15_13_port, A2 => n27026, ZN => 
                           N548);
   U2654 : AND2_X1 port map( A1 => regs_nxt_15_14_port, A2 => n26989, ZN => 
                           N549);
   U2655 : AND2_X1 port map( A1 => regs_nxt_15_15_port, A2 => n26985, ZN => 
                           N550);
   U2656 : AND2_X1 port map( A1 => regs_nxt_15_16_port, A2 => n26981, ZN => 
                           N551);
   U2657 : AND2_X1 port map( A1 => regs_nxt_15_17_port, A2 => n26981, ZN => 
                           N552);
   U2658 : AND2_X1 port map( A1 => regs_nxt_15_18_port, A2 => n26981, ZN => 
                           N553);
   U2659 : AND2_X1 port map( A1 => regs_nxt_15_19_port, A2 => n26981, ZN => 
                           N554);
   U2660 : AND2_X1 port map( A1 => regs_nxt_15_20_port, A2 => n26981, ZN => 
                           N555);
   U2661 : AND2_X1 port map( A1 => regs_nxt_15_21_port, A2 => n26981, ZN => 
                           N556);
   U2662 : AND2_X1 port map( A1 => regs_nxt_15_22_port, A2 => n26981, ZN => 
                           N557);
   U2663 : AND2_X1 port map( A1 => regs_nxt_15_23_port, A2 => n26981, ZN => 
                           N558);
   U2664 : AND2_X1 port map( A1 => regs_nxt_15_24_port, A2 => n26981, ZN => 
                           N559);
   U2665 : AND2_X1 port map( A1 => regs_nxt_15_25_port, A2 => n26981, ZN => 
                           N560);
   U2666 : AND2_X1 port map( A1 => regs_nxt_15_26_port, A2 => n26982, ZN => 
                           N561);
   U2667 : AND2_X1 port map( A1 => regs_nxt_15_27_port, A2 => n26982, ZN => 
                           N562);
   U2668 : AND2_X1 port map( A1 => regs_nxt_15_28_port, A2 => n26982, ZN => 
                           N563);
   U2669 : AND2_X1 port map( A1 => regs_nxt_15_29_port, A2 => n26982, ZN => 
                           N564);
   U2670 : AND2_X1 port map( A1 => regs_nxt_15_30_port, A2 => n26982, ZN => 
                           N565);
   U2671 : AND2_X1 port map( A1 => regs_nxt_15_31_port, A2 => n26982, ZN => 
                           N566);
   U2672 : AND2_X1 port map( A1 => regs_nxt_14_0_port, A2 => n26982, ZN => N567
                           );
   U2673 : AND2_X1 port map( A1 => regs_nxt_14_1_port, A2 => n26982, ZN => N568
                           );
   U2674 : AND2_X1 port map( A1 => regs_nxt_14_2_port, A2 => n26982, ZN => N569
                           );
   U2675 : AND2_X1 port map( A1 => regs_nxt_14_3_port, A2 => n26982, ZN => N570
                           );
   U2676 : AND2_X1 port map( A1 => regs_nxt_14_4_port, A2 => n26982, ZN => N571
                           );
   U2677 : AND2_X1 port map( A1 => regs_nxt_14_5_port, A2 => n26982, ZN => N572
                           );
   U2678 : AND2_X1 port map( A1 => regs_nxt_14_6_port, A2 => n26982, ZN => N573
                           );
   U2679 : AND2_X1 port map( A1 => regs_nxt_14_7_port, A2 => n26982, ZN => N574
                           );
   U2680 : AND2_X1 port map( A1 => regs_nxt_14_8_port, A2 => n26982, ZN => N575
                           );
   U2681 : AND2_X1 port map( A1 => regs_nxt_14_9_port, A2 => n26982, ZN => N576
                           );
   U2682 : AND2_X1 port map( A1 => regs_nxt_14_10_port, A2 => n26982, ZN => 
                           N577);
   U2683 : AND2_X1 port map( A1 => regs_nxt_14_11_port, A2 => n26983, ZN => 
                           N578);
   U2684 : AND2_X1 port map( A1 => regs_nxt_14_12_port, A2 => n26983, ZN => 
                           N579);
   U2685 : AND2_X1 port map( A1 => regs_nxt_14_13_port, A2 => n26983, ZN => 
                           N580);
   U2686 : AND2_X1 port map( A1 => regs_nxt_14_14_port, A2 => n26983, ZN => 
                           N581);
   U2687 : AND2_X1 port map( A1 => regs_nxt_14_15_port, A2 => n26983, ZN => 
                           N582);
   U2688 : AND2_X1 port map( A1 => regs_nxt_14_16_port, A2 => n26983, ZN => 
                           N583);
   U2689 : AND2_X1 port map( A1 => regs_nxt_14_17_port, A2 => n26983, ZN => 
                           N584);
   U2690 : AND2_X1 port map( A1 => regs_nxt_14_18_port, A2 => n26983, ZN => 
                           N585);
   U2691 : AND2_X1 port map( A1 => regs_nxt_14_19_port, A2 => n26983, ZN => 
                           N586);
   U2692 : AND2_X1 port map( A1 => regs_nxt_14_20_port, A2 => n26983, ZN => 
                           N587);
   U2693 : AND2_X1 port map( A1 => regs_nxt_14_21_port, A2 => n26983, ZN => 
                           N588);
   U2694 : AND2_X1 port map( A1 => regs_nxt_14_22_port, A2 => n26983, ZN => 
                           N589);
   U2695 : AND2_X1 port map( A1 => regs_nxt_14_23_port, A2 => n26983, ZN => 
                           N590);
   U2696 : AND2_X1 port map( A1 => regs_nxt_14_24_port, A2 => n26983, ZN => 
                           N591);
   U2697 : AND2_X1 port map( A1 => regs_nxt_14_25_port, A2 => n26983, ZN => 
                           N592);
   U2698 : AND2_X1 port map( A1 => regs_nxt_14_26_port, A2 => n26983, ZN => 
                           N593);
   U2699 : AND2_X1 port map( A1 => regs_nxt_14_27_port, A2 => n26984, ZN => 
                           N594);
   U2700 : AND2_X1 port map( A1 => regs_nxt_14_28_port, A2 => n26984, ZN => 
                           N595);
   U2701 : AND2_X1 port map( A1 => regs_nxt_14_29_port, A2 => n26984, ZN => 
                           N596);
   U2702 : AND2_X1 port map( A1 => regs_nxt_14_30_port, A2 => n26984, ZN => 
                           N597);
   U2703 : AND2_X1 port map( A1 => regs_nxt_14_31_port, A2 => n26984, ZN => 
                           N598);
   U2704 : AND2_X1 port map( A1 => regs_nxt_13_0_port, A2 => n26984, ZN => N599
                           );
   U2705 : AND2_X1 port map( A1 => regs_nxt_13_1_port, A2 => n26984, ZN => N600
                           );
   U2706 : AND2_X1 port map( A1 => regs_nxt_13_2_port, A2 => n26984, ZN => N601
                           );
   U2707 : AND2_X1 port map( A1 => regs_nxt_13_3_port, A2 => n26984, ZN => N602
                           );
   U2708 : AND2_X1 port map( A1 => regs_nxt_13_4_port, A2 => n26984, ZN => N603
                           );
   U2709 : AND2_X1 port map( A1 => regs_nxt_13_5_port, A2 => n26984, ZN => N604
                           );
   U2710 : AND2_X1 port map( A1 => regs_nxt_13_6_port, A2 => n26984, ZN => N605
                           );
   U2711 : AND2_X1 port map( A1 => regs_nxt_13_7_port, A2 => n26984, ZN => N606
                           );
   U2712 : AND2_X1 port map( A1 => regs_nxt_13_8_port, A2 => n26984, ZN => N607
                           );
   U2713 : AND2_X1 port map( A1 => regs_nxt_13_9_port, A2 => n26984, ZN => N608
                           );
   U2714 : AND2_X1 port map( A1 => regs_nxt_13_10_port, A2 => n26984, ZN => 
                           N609);
   U2715 : AND2_X1 port map( A1 => regs_nxt_13_11_port, A2 => n26985, ZN => 
                           N610);
   U2716 : AND2_X1 port map( A1 => regs_nxt_13_12_port, A2 => n26985, ZN => 
                           N611);
   U2717 : AND2_X1 port map( A1 => regs_nxt_13_13_port, A2 => n26985, ZN => 
                           N612);
   U2718 : AND2_X1 port map( A1 => regs_nxt_13_14_port, A2 => n26985, ZN => 
                           N613);
   U2719 : AND2_X1 port map( A1 => regs_nxt_13_15_port, A2 => n26985, ZN => 
                           N614);
   U2720 : AND2_X1 port map( A1 => regs_nxt_13_16_port, A2 => n26985, ZN => 
                           N615);
   U2721 : AND2_X1 port map( A1 => regs_nxt_13_17_port, A2 => n26985, ZN => 
                           N616);
   U2722 : AND2_X1 port map( A1 => regs_nxt_13_18_port, A2 => n26985, ZN => 
                           N617);
   U2723 : AND2_X1 port map( A1 => regs_nxt_13_19_port, A2 => n26985, ZN => 
                           N618);
   U2724 : AND2_X1 port map( A1 => regs_nxt_13_20_port, A2 => n26985, ZN => 
                           N619);
   U2725 : AND2_X1 port map( A1 => regs_nxt_13_21_port, A2 => n26985, ZN => 
                           N620);
   U2726 : AND2_X1 port map( A1 => regs_nxt_13_22_port, A2 => n26985, ZN => 
                           N621);
   U2727 : AND2_X1 port map( A1 => regs_nxt_13_23_port, A2 => n26985, ZN => 
                           N622);
   U2728 : AND2_X1 port map( A1 => regs_nxt_13_24_port, A2 => n26985, ZN => 
                           N623);
   U2729 : AND2_X1 port map( A1 => regs_nxt_13_25_port, A2 => n26985, ZN => 
                           N624);
   U2730 : AND2_X1 port map( A1 => regs_nxt_13_26_port, A2 => n26985, ZN => 
                           N625);
   U2731 : AND2_X1 port map( A1 => regs_nxt_13_27_port, A2 => n26986, ZN => 
                           N626);
   U2732 : AND2_X1 port map( A1 => regs_nxt_13_28_port, A2 => n26986, ZN => 
                           N627);
   U2733 : AND2_X1 port map( A1 => regs_nxt_13_29_port, A2 => n26986, ZN => 
                           N628);
   U2734 : AND2_X1 port map( A1 => regs_nxt_13_30_port, A2 => n26986, ZN => 
                           N629);
   U2735 : AND2_X1 port map( A1 => regs_nxt_13_31_port, A2 => n26986, ZN => 
                           N630);
   U2736 : AND2_X1 port map( A1 => regs_nxt_12_0_port, A2 => n26986, ZN => N631
                           );
   U2737 : AND2_X1 port map( A1 => regs_nxt_12_1_port, A2 => n26986, ZN => N632
                           );
   U2738 : AND2_X1 port map( A1 => regs_nxt_12_2_port, A2 => n26986, ZN => N633
                           );
   U2739 : AND2_X1 port map( A1 => regs_nxt_12_3_port, A2 => n26986, ZN => N634
                           );
   U2740 : AND2_X1 port map( A1 => regs_nxt_12_4_port, A2 => n26986, ZN => N635
                           );
   U2741 : AND2_X1 port map( A1 => regs_nxt_12_5_port, A2 => n26986, ZN => N636
                           );
   U2742 : AND2_X1 port map( A1 => regs_nxt_12_6_port, A2 => n26986, ZN => N637
                           );
   U2743 : AND2_X1 port map( A1 => regs_nxt_12_7_port, A2 => n26986, ZN => N638
                           );
   U2744 : AND2_X1 port map( A1 => regs_nxt_12_8_port, A2 => n26986, ZN => N639
                           );
   U2745 : AND2_X1 port map( A1 => regs_nxt_12_9_port, A2 => n26986, ZN => N640
                           );
   U2746 : AND2_X1 port map( A1 => regs_nxt_12_10_port, A2 => n26986, ZN => 
                           N641);
   U2747 : AND2_X1 port map( A1 => regs_nxt_12_11_port, A2 => n26987, ZN => 
                           N642);
   U2748 : AND2_X1 port map( A1 => regs_nxt_12_12_port, A2 => n26987, ZN => 
                           N643);
   U2749 : AND2_X1 port map( A1 => regs_nxt_12_13_port, A2 => n26987, ZN => 
                           N644);
   U2750 : AND2_X1 port map( A1 => regs_nxt_12_14_port, A2 => n26987, ZN => 
                           N645);
   U2751 : AND2_X1 port map( A1 => regs_nxt_12_15_port, A2 => n26987, ZN => 
                           N646);
   U2752 : AND2_X1 port map( A1 => regs_nxt_12_16_port, A2 => n26987, ZN => 
                           N647);
   U2753 : AND2_X1 port map( A1 => regs_nxt_12_17_port, A2 => n26987, ZN => 
                           N648);
   U2754 : AND2_X1 port map( A1 => regs_nxt_12_18_port, A2 => n26987, ZN => 
                           N649);
   U2755 : AND2_X1 port map( A1 => regs_nxt_12_19_port, A2 => n26987, ZN => 
                           N650);
   U2756 : AND2_X1 port map( A1 => regs_nxt_12_20_port, A2 => n26987, ZN => 
                           N651);
   U2757 : AND2_X1 port map( A1 => regs_nxt_12_21_port, A2 => n26987, ZN => 
                           N652);
   U2758 : AND2_X1 port map( A1 => regs_nxt_12_22_port, A2 => n26987, ZN => 
                           N653);
   U2759 : AND2_X1 port map( A1 => regs_nxt_12_23_port, A2 => n26987, ZN => 
                           N654);
   U2760 : AND2_X1 port map( A1 => regs_nxt_12_24_port, A2 => n26987, ZN => 
                           N655);
   U2761 : AND2_X1 port map( A1 => regs_nxt_12_25_port, A2 => n26987, ZN => 
                           N656);
   U2762 : AND2_X1 port map( A1 => regs_nxt_12_26_port, A2 => n26987, ZN => 
                           N657);
   U2763 : AND2_X1 port map( A1 => regs_nxt_12_27_port, A2 => n26987, ZN => 
                           N658);
   U2764 : AND2_X1 port map( A1 => regs_nxt_12_28_port, A2 => n26988, ZN => 
                           N659);
   U2765 : AND2_X1 port map( A1 => regs_nxt_12_29_port, A2 => n26988, ZN => 
                           N660);
   U2766 : AND2_X1 port map( A1 => regs_nxt_12_30_port, A2 => n26988, ZN => 
                           N661);
   U2767 : AND2_X1 port map( A1 => regs_nxt_12_31_port, A2 => n26988, ZN => 
                           N662);
   U2768 : AND2_X1 port map( A1 => regs_nxt_11_0_port, A2 => n26988, ZN => N663
                           );
   U2769 : AND2_X1 port map( A1 => regs_nxt_11_1_port, A2 => n26988, ZN => N664
                           );
   U2770 : AND2_X1 port map( A1 => regs_nxt_11_2_port, A2 => n26988, ZN => N665
                           );
   U2771 : AND2_X1 port map( A1 => regs_nxt_11_3_port, A2 => n26988, ZN => N666
                           );
   U2772 : AND2_X1 port map( A1 => regs_nxt_11_4_port, A2 => n26988, ZN => N667
                           );
   U2773 : AND2_X1 port map( A1 => regs_nxt_11_5_port, A2 => n26988, ZN => N668
                           );
   U2774 : AND2_X1 port map( A1 => regs_nxt_11_6_port, A2 => n26988, ZN => N669
                           );
   U2775 : AND2_X1 port map( A1 => regs_nxt_11_7_port, A2 => n26988, ZN => N670
                           );
   U2776 : AND2_X1 port map( A1 => regs_nxt_11_8_port, A2 => n26988, ZN => N671
                           );
   U2777 : AND2_X1 port map( A1 => regs_nxt_11_9_port, A2 => n26988, ZN => N672
                           );
   U2778 : AND2_X1 port map( A1 => regs_nxt_11_10_port, A2 => n26988, ZN => 
                           N673);
   U2779 : AND2_X1 port map( A1 => regs_nxt_11_11_port, A2 => n26988, ZN => 
                           N674);
   U2780 : AND2_X1 port map( A1 => regs_nxt_11_12_port, A2 => n26989, ZN => 
                           N675);
   U2781 : AND2_X1 port map( A1 => regs_nxt_11_13_port, A2 => n26989, ZN => 
                           N676);
   U2782 : AND2_X1 port map( A1 => regs_nxt_11_14_port, A2 => n26989, ZN => 
                           N677);
   U2783 : AND2_X1 port map( A1 => regs_nxt_11_15_port, A2 => n26989, ZN => 
                           N678);
   U2784 : AND2_X1 port map( A1 => regs_nxt_11_16_port, A2 => n26989, ZN => 
                           N679);
   U2785 : AND2_X1 port map( A1 => regs_nxt_11_17_port, A2 => n26989, ZN => 
                           N680);
   U2786 : AND2_X1 port map( A1 => regs_nxt_11_18_port, A2 => n26989, ZN => 
                           N681);
   U2787 : AND2_X1 port map( A1 => regs_nxt_11_19_port, A2 => n26989, ZN => 
                           N682);
   U2788 : AND2_X1 port map( A1 => regs_nxt_11_20_port, A2 => n26977, ZN => 
                           N683);
   U2789 : AND2_X1 port map( A1 => regs_nxt_11_21_port, A2 => n26975, ZN => 
                           N684);
   U2790 : AND2_X1 port map( A1 => regs_nxt_11_22_port, A2 => n26976, ZN => 
                           N685);
   U2791 : AND2_X1 port map( A1 => regs_nxt_11_23_port, A2 => n26974, ZN => 
                           N686);
   U2792 : AND2_X1 port map( A1 => regs_nxt_11_24_port, A2 => n26976, ZN => 
                           N687);
   U2793 : AND2_X1 port map( A1 => regs_nxt_11_25_port, A2 => n26975, ZN => 
                           N688);
   U2794 : AND2_X1 port map( A1 => regs_nxt_11_26_port, A2 => n26975, ZN => 
                           N689);
   U2795 : AND2_X1 port map( A1 => regs_nxt_11_27_port, A2 => n26975, ZN => 
                           N690);
   U2796 : AND2_X1 port map( A1 => regs_nxt_11_28_port, A2 => n26975, ZN => 
                           N691);
   U2797 : AND2_X1 port map( A1 => regs_nxt_11_29_port, A2 => n26975, ZN => 
                           N692);
   U2798 : AND2_X1 port map( A1 => regs_nxt_11_30_port, A2 => n26975, ZN => 
                           N693);
   U2799 : AND2_X1 port map( A1 => regs_nxt_11_31_port, A2 => n26975, ZN => 
                           N694);
   U2800 : AND2_X1 port map( A1 => regs_nxt_10_0_port, A2 => n26975, ZN => N695
                           );
   U2801 : AND2_X1 port map( A1 => regs_nxt_10_1_port, A2 => n26975, ZN => N696
                           );
   U2802 : AND2_X1 port map( A1 => regs_nxt_10_2_port, A2 => n26975, ZN => N697
                           );
   U2803 : AND2_X1 port map( A1 => regs_nxt_10_3_port, A2 => n26975, ZN => N698
                           );
   U2804 : AND2_X1 port map( A1 => regs_nxt_10_4_port, A2 => n26976, ZN => N699
                           );
   U2805 : AND2_X1 port map( A1 => regs_nxt_10_5_port, A2 => n26975, ZN => N700
                           );
   U2806 : AND2_X1 port map( A1 => regs_nxt_10_6_port, A2 => n26975, ZN => N701
                           );
   U2807 : AND2_X1 port map( A1 => regs_nxt_10_7_port, A2 => n26975, ZN => N702
                           );
   U2808 : AND2_X1 port map( A1 => regs_nxt_10_8_port, A2 => n26976, ZN => N703
                           );
   U2809 : AND2_X1 port map( A1 => regs_nxt_10_9_port, A2 => n26975, ZN => N704
                           );
   U2810 : AND2_X1 port map( A1 => regs_nxt_10_10_port, A2 => n26976, ZN => 
                           N705);
   U2811 : AND2_X1 port map( A1 => regs_nxt_10_11_port, A2 => n26976, ZN => 
                           N706);
   U2812 : AND2_X1 port map( A1 => regs_nxt_10_12_port, A2 => n26976, ZN => 
                           N707);
   U2813 : AND2_X1 port map( A1 => regs_nxt_10_13_port, A2 => n26976, ZN => 
                           N708);
   U2814 : AND2_X1 port map( A1 => regs_nxt_10_14_port, A2 => n26976, ZN => 
                           N709);
   U2815 : AND2_X1 port map( A1 => regs_nxt_10_15_port, A2 => n26976, ZN => 
                           N710);
   U2816 : AND2_X1 port map( A1 => regs_nxt_10_16_port, A2 => n26976, ZN => 
                           N711);
   U2817 : AND2_X1 port map( A1 => regs_nxt_10_17_port, A2 => n26976, ZN => 
                           N712);
   U2818 : AND2_X1 port map( A1 => regs_nxt_10_18_port, A2 => n26976, ZN => 
                           N713);
   U2819 : AND2_X1 port map( A1 => regs_nxt_10_19_port, A2 => n26976, ZN => 
                           N714);
   U2820 : AND2_X1 port map( A1 => regs_nxt_10_20_port, A2 => n26976, ZN => 
                           N715);
   U2821 : AND2_X1 port map( A1 => regs_nxt_10_21_port, A2 => n26976, ZN => 
                           N716);
   U2822 : AND2_X1 port map( A1 => regs_nxt_10_22_port, A2 => n26977, ZN => 
                           N717);
   U2823 : AND2_X1 port map( A1 => regs_nxt_10_23_port, A2 => n26976, ZN => 
                           N718);
   U2824 : AND2_X1 port map( A1 => regs_nxt_10_24_port, A2 => n26977, ZN => 
                           N719);
   U2825 : AND2_X1 port map( A1 => regs_nxt_10_25_port, A2 => n26977, ZN => 
                           N720);
   U2826 : AND2_X1 port map( A1 => regs_nxt_10_26_port, A2 => n26977, ZN => 
                           N721);
   U2827 : AND2_X1 port map( A1 => regs_nxt_10_27_port, A2 => n26977, ZN => 
                           N722);
   U2828 : AND2_X1 port map( A1 => regs_nxt_10_28_port, A2 => n26977, ZN => 
                           N723);
   U2829 : AND2_X1 port map( A1 => regs_nxt_10_29_port, A2 => n26977, ZN => 
                           N724);
   U2830 : AND2_X1 port map( A1 => regs_nxt_10_30_port, A2 => n26977, ZN => 
                           N725);
   U2831 : AND2_X1 port map( A1 => regs_nxt_10_31_port, A2 => n26977, ZN => 
                           N726);
   U2832 : AND2_X1 port map( A1 => regs_nxt_9_0_port, A2 => n26977, ZN => N727)
                           ;
   U2833 : AND2_X1 port map( A1 => regs_nxt_9_1_port, A2 => n26977, ZN => N728)
                           ;
   U2834 : AND2_X1 port map( A1 => regs_nxt_9_2_port, A2 => n26977, ZN => N729)
                           ;
   U2835 : AND2_X1 port map( A1 => regs_nxt_9_3_port, A2 => n26977, ZN => N730)
                           ;
   U2836 : AND2_X1 port map( A1 => regs_nxt_9_4_port, A2 => n26977, ZN => N731)
                           ;
   U2837 : AND2_X1 port map( A1 => regs_nxt_9_5_port, A2 => n26977, ZN => N732)
                           ;
   U2838 : AND2_X1 port map( A1 => regs_nxt_9_6_port, A2 => n26978, ZN => N733)
                           ;
   U2839 : AND2_X1 port map( A1 => regs_nxt_9_7_port, A2 => n26978, ZN => N734)
                           ;
   U2840 : AND2_X1 port map( A1 => regs_nxt_9_8_port, A2 => n26978, ZN => N735)
                           ;
   U2841 : AND2_X1 port map( A1 => regs_nxt_9_9_port, A2 => n26978, ZN => N736)
                           ;
   U2842 : AND2_X1 port map( A1 => regs_nxt_9_10_port, A2 => n26978, ZN => N737
                           );
   U2843 : AND2_X1 port map( A1 => regs_nxt_9_11_port, A2 => n26978, ZN => N738
                           );
   U2844 : AND2_X1 port map( A1 => regs_nxt_9_12_port, A2 => n26978, ZN => N739
                           );
   U2845 : AND2_X1 port map( A1 => regs_nxt_9_13_port, A2 => n26978, ZN => N740
                           );
   U2846 : AND2_X1 port map( A1 => regs_nxt_9_14_port, A2 => n26978, ZN => N741
                           );
   U2847 : AND2_X1 port map( A1 => regs_nxt_9_15_port, A2 => n26978, ZN => N742
                           );
   U2848 : AND2_X1 port map( A1 => regs_nxt_9_16_port, A2 => n26978, ZN => N743
                           );
   U2849 : AND2_X1 port map( A1 => regs_nxt_9_17_port, A2 => n26978, ZN => N744
                           );
   U2850 : AND2_X1 port map( A1 => regs_nxt_9_18_port, A2 => n26978, ZN => N745
                           );
   U2851 : AND2_X1 port map( A1 => regs_nxt_9_19_port, A2 => n26978, ZN => N746
                           );
   U2852 : AND2_X1 port map( A1 => regs_nxt_9_20_port, A2 => n26978, ZN => N747
                           );
   U2853 : AND2_X1 port map( A1 => regs_nxt_9_21_port, A2 => n26978, ZN => N748
                           );
   U2854 : AND2_X1 port map( A1 => regs_nxt_9_22_port, A2 => n26978, ZN => N749
                           );
   U2855 : AND2_X1 port map( A1 => regs_nxt_9_23_port, A2 => n26979, ZN => N750
                           );
   U2856 : AND2_X1 port map( A1 => regs_nxt_9_24_port, A2 => n26979, ZN => N751
                           );
   U2857 : AND2_X1 port map( A1 => regs_nxt_9_25_port, A2 => n26979, ZN => N752
                           );
   U2858 : AND2_X1 port map( A1 => regs_nxt_9_26_port, A2 => n26979, ZN => N753
                           );
   U2859 : AND2_X1 port map( A1 => regs_nxt_9_27_port, A2 => n26979, ZN => N754
                           );
   U2860 : AND2_X1 port map( A1 => regs_nxt_9_28_port, A2 => n26979, ZN => N755
                           );
   U2861 : AND2_X1 port map( A1 => regs_nxt_9_29_port, A2 => n26979, ZN => N756
                           );
   U2862 : AND2_X1 port map( A1 => regs_nxt_9_30_port, A2 => n26979, ZN => N757
                           );
   U2863 : AND2_X1 port map( A1 => regs_nxt_9_31_port, A2 => n26979, ZN => N758
                           );
   U2864 : AND2_X1 port map( A1 => regs_nxt_8_0_port, A2 => n26979, ZN => N759)
                           ;
   U2865 : AND2_X1 port map( A1 => regs_nxt_8_1_port, A2 => n26979, ZN => N760)
                           ;
   U2866 : AND2_X1 port map( A1 => regs_nxt_8_2_port, A2 => n26979, ZN => N761)
                           ;
   U2867 : AND2_X1 port map( A1 => regs_nxt_8_3_port, A2 => n26979, ZN => N762)
                           ;
   U2868 : AND2_X1 port map( A1 => regs_nxt_8_4_port, A2 => n26979, ZN => N763)
                           ;
   U2869 : AND2_X1 port map( A1 => regs_nxt_8_5_port, A2 => n26979, ZN => N764)
                           ;
   U2870 : AND2_X1 port map( A1 => regs_nxt_8_6_port, A2 => n26979, ZN => N765)
                           ;
   U2871 : AND2_X1 port map( A1 => regs_nxt_8_7_port, A2 => n26980, ZN => N766)
                           ;
   U2872 : AND2_X1 port map( A1 => regs_nxt_8_8_port, A2 => n26980, ZN => N767)
                           ;
   U2873 : AND2_X1 port map( A1 => regs_nxt_8_9_port, A2 => n26980, ZN => N768)
                           ;
   U2874 : AND2_X1 port map( A1 => regs_nxt_8_10_port, A2 => n26980, ZN => N769
                           );
   U2875 : AND2_X1 port map( A1 => regs_nxt_8_11_port, A2 => n26980, ZN => N770
                           );
   U2876 : AND2_X1 port map( A1 => regs_nxt_8_12_port, A2 => n26980, ZN => N771
                           );
   U2877 : AND2_X1 port map( A1 => regs_nxt_8_13_port, A2 => n26980, ZN => N772
                           );
   U2878 : AND2_X1 port map( A1 => regs_nxt_8_14_port, A2 => n26980, ZN => N773
                           );
   U2879 : AND2_X1 port map( A1 => regs_nxt_8_15_port, A2 => n26980, ZN => N774
                           );
   U2880 : AND2_X1 port map( A1 => regs_nxt_8_16_port, A2 => n26980, ZN => N775
                           );
   U2881 : AND2_X1 port map( A1 => regs_nxt_8_17_port, A2 => n26980, ZN => N776
                           );
   U2882 : AND2_X1 port map( A1 => regs_nxt_8_18_port, A2 => n26980, ZN => N777
                           );
   U2883 : AND2_X1 port map( A1 => regs_nxt_8_19_port, A2 => n26980, ZN => N778
                           );
   U2884 : AND2_X1 port map( A1 => regs_nxt_8_20_port, A2 => n26980, ZN => N779
                           );
   U2885 : AND2_X1 port map( A1 => regs_nxt_8_21_port, A2 => n26980, ZN => N780
                           );
   U2886 : AND2_X1 port map( A1 => regs_nxt_8_22_port, A2 => n26980, ZN => N781
                           );
   U2887 : AND2_X1 port map( A1 => regs_nxt_8_23_port, A2 => n26981, ZN => N782
                           );
   U2888 : AND2_X1 port map( A1 => regs_nxt_8_24_port, A2 => n26981, ZN => N783
                           );
   U2889 : AND2_X1 port map( A1 => regs_nxt_8_25_port, A2 => n26981, ZN => N784
                           );
   U2890 : AND2_X1 port map( A1 => regs_nxt_8_26_port, A2 => n26981, ZN => N785
                           );
   U2891 : AND2_X1 port map( A1 => regs_nxt_8_27_port, A2 => n26981, ZN => N786
                           );
   U2892 : AND2_X1 port map( A1 => regs_nxt_8_28_port, A2 => n26981, ZN => N787
                           );
   U2893 : AND2_X1 port map( A1 => regs_nxt_8_29_port, A2 => n27000, ZN => N788
                           );
   U2894 : AND2_X1 port map( A1 => regs_nxt_8_30_port, A2 => n26996, ZN => N789
                           );
   U2895 : AND2_X1 port map( A1 => regs_nxt_8_31_port, A2 => n26997, ZN => N790
                           );
   U2896 : AND2_X1 port map( A1 => regs_nxt_7_0_port, A2 => n26997, ZN => N791)
                           ;
   U2897 : AND2_X1 port map( A1 => regs_nxt_7_1_port, A2 => n26997, ZN => N792)
                           ;
   U2898 : AND2_X1 port map( A1 => regs_nxt_7_2_port, A2 => n26997, ZN => N793)
                           ;
   U2899 : AND2_X1 port map( A1 => regs_nxt_7_3_port, A2 => n26997, ZN => N794)
                           ;
   U2900 : AND2_X1 port map( A1 => regs_nxt_7_4_port, A2 => n26997, ZN => N795)
                           ;
   U2901 : AND2_X1 port map( A1 => regs_nxt_7_5_port, A2 => n26997, ZN => N796)
                           ;
   U2902 : AND2_X1 port map( A1 => regs_nxt_7_6_port, A2 => n26997, ZN => N797)
                           ;
   U2903 : AND2_X1 port map( A1 => regs_nxt_7_7_port, A2 => n26997, ZN => N798)
                           ;
   U2904 : AND2_X1 port map( A1 => regs_nxt_7_8_port, A2 => n26997, ZN => N799)
                           ;
   U2905 : AND2_X1 port map( A1 => regs_nxt_7_9_port, A2 => n26997, ZN => N800)
                           ;
   U2906 : AND2_X1 port map( A1 => regs_nxt_7_10_port, A2 => n26997, ZN => N801
                           );
   U2907 : AND2_X1 port map( A1 => regs_nxt_7_11_port, A2 => n26997, ZN => N802
                           );
   U2908 : AND2_X1 port map( A1 => regs_nxt_7_12_port, A2 => n26997, ZN => N803
                           );
   U2909 : AND2_X1 port map( A1 => regs_nxt_7_13_port, A2 => n26997, ZN => N804
                           );
   U2910 : AND2_X1 port map( A1 => regs_nxt_7_14_port, A2 => n26997, ZN => N805
                           );
   U2911 : AND2_X1 port map( A1 => regs_nxt_7_15_port, A2 => n26997, ZN => N806
                           );
   U2912 : AND2_X1 port map( A1 => regs_nxt_7_16_port, A2 => n26998, ZN => N807
                           );
   U2913 : AND2_X1 port map( A1 => regs_nxt_7_17_port, A2 => n26998, ZN => N808
                           );
   U2914 : AND2_X1 port map( A1 => regs_nxt_7_18_port, A2 => n26998, ZN => N809
                           );
   U2915 : AND2_X1 port map( A1 => regs_nxt_7_19_port, A2 => n26998, ZN => N810
                           );
   U2916 : AND2_X1 port map( A1 => regs_nxt_7_20_port, A2 => n26998, ZN => N811
                           );
   U2917 : AND2_X1 port map( A1 => regs_nxt_7_21_port, A2 => n26998, ZN => N812
                           );
   U2918 : AND2_X1 port map( A1 => regs_nxt_7_22_port, A2 => n26998, ZN => N813
                           );
   U2919 : AND2_X1 port map( A1 => regs_nxt_7_23_port, A2 => n26998, ZN => N814
                           );
   U2920 : AND2_X1 port map( A1 => regs_nxt_7_24_port, A2 => n26998, ZN => N815
                           );
   U2921 : AND2_X1 port map( A1 => regs_nxt_7_25_port, A2 => n26998, ZN => N816
                           );
   U2922 : AND2_X1 port map( A1 => regs_nxt_7_26_port, A2 => n26998, ZN => N817
                           );
   U2923 : AND2_X1 port map( A1 => regs_nxt_7_27_port, A2 => n26998, ZN => N818
                           );
   U2924 : AND2_X1 port map( A1 => regs_nxt_7_28_port, A2 => n26998, ZN => N819
                           );
   U2925 : AND2_X1 port map( A1 => regs_nxt_7_29_port, A2 => n26998, ZN => N820
                           );
   U2926 : AND2_X1 port map( A1 => regs_nxt_7_30_port, A2 => n26998, ZN => N821
                           );
   U2927 : AND2_X1 port map( A1 => regs_nxt_7_31_port, A2 => n26998, ZN => N822
                           );
   U2928 : AND2_X1 port map( A1 => regs_nxt_6_0_port, A2 => n26999, ZN => N823)
                           ;
   U2929 : AND2_X1 port map( A1 => regs_nxt_6_1_port, A2 => n26999, ZN => N824)
                           ;
   U2930 : AND2_X1 port map( A1 => regs_nxt_6_2_port, A2 => n26999, ZN => N825)
                           ;
   U2931 : AND2_X1 port map( A1 => regs_nxt_6_3_port, A2 => n26999, ZN => N826)
                           ;
   U2932 : AND2_X1 port map( A1 => regs_nxt_6_4_port, A2 => n26999, ZN => N827)
                           ;
   U2933 : AND2_X1 port map( A1 => regs_nxt_6_5_port, A2 => n26999, ZN => N828)
                           ;
   U2934 : AND2_X1 port map( A1 => regs_nxt_6_6_port, A2 => n26999, ZN => N829)
                           ;
   U2935 : AND2_X1 port map( A1 => regs_nxt_6_7_port, A2 => n26999, ZN => N830)
                           ;
   U2936 : AND2_X1 port map( A1 => regs_nxt_6_8_port, A2 => n26999, ZN => N831)
                           ;
   U2937 : AND2_X1 port map( A1 => regs_nxt_6_9_port, A2 => n26999, ZN => N832)
                           ;
   U2938 : AND2_X1 port map( A1 => regs_nxt_6_10_port, A2 => n26999, ZN => N833
                           );
   U2939 : AND2_X1 port map( A1 => regs_nxt_6_11_port, A2 => n26999, ZN => N834
                           );
   U2940 : AND2_X1 port map( A1 => regs_nxt_6_12_port, A2 => n26999, ZN => N835
                           );
   U2941 : AND2_X1 port map( A1 => regs_nxt_6_13_port, A2 => n26999, ZN => N836
                           );
   U2942 : AND2_X1 port map( A1 => regs_nxt_6_14_port, A2 => n26999, ZN => N837
                           );
   U2943 : AND2_X1 port map( A1 => regs_nxt_6_15_port, A2 => n26999, ZN => N838
                           );
   U2944 : AND2_X1 port map( A1 => regs_nxt_6_16_port, A2 => n26999, ZN => N839
                           );
   U2945 : AND2_X1 port map( A1 => regs_nxt_6_17_port, A2 => n27000, ZN => N840
                           );
   U2946 : AND2_X1 port map( A1 => regs_nxt_6_18_port, A2 => n27000, ZN => N841
                           );
   U2947 : AND2_X1 port map( A1 => regs_nxt_6_19_port, A2 => n27000, ZN => N842
                           );
   U2948 : AND2_X1 port map( A1 => regs_nxt_6_20_port, A2 => n27000, ZN => N843
                           );
   U2949 : AND2_X1 port map( A1 => regs_nxt_6_21_port, A2 => n27000, ZN => N844
                           );
   U2950 : AND2_X1 port map( A1 => regs_nxt_6_22_port, A2 => n27000, ZN => N845
                           );
   U2951 : AND2_X1 port map( A1 => regs_nxt_6_23_port, A2 => n27000, ZN => N846
                           );
   U2952 : AND2_X1 port map( A1 => regs_nxt_6_24_port, A2 => n27000, ZN => N847
                           );
   U2953 : AND2_X1 port map( A1 => regs_nxt_6_25_port, A2 => n27000, ZN => N848
                           );
   U2954 : AND2_X1 port map( A1 => regs_nxt_6_26_port, A2 => n27000, ZN => N849
                           );
   U2955 : AND2_X1 port map( A1 => regs_nxt_6_27_port, A2 => n27000, ZN => N850
                           );
   U2956 : AND2_X1 port map( A1 => regs_nxt_6_28_port, A2 => n27000, ZN => N851
                           );
   U2957 : AND2_X1 port map( A1 => regs_nxt_6_29_port, A2 => n27000, ZN => N852
                           );
   U2958 : AND2_X1 port map( A1 => regs_nxt_6_30_port, A2 => n27000, ZN => N853
                           );
   U2959 : AND2_X1 port map( A1 => regs_nxt_6_31_port, A2 => n27000, ZN => N854
                           );
   U2960 : AND2_X1 port map( A1 => regs_nxt_5_0_port, A2 => n27001, ZN => N855)
                           ;
   U2961 : AND2_X1 port map( A1 => regs_nxt_5_1_port, A2 => n27001, ZN => N856)
                           ;
   U2962 : AND2_X1 port map( A1 => regs_nxt_5_2_port, A2 => n27001, ZN => N857)
                           ;
   U2963 : AND2_X1 port map( A1 => regs_nxt_5_3_port, A2 => n27001, ZN => N858)
                           ;
   U2964 : AND2_X1 port map( A1 => regs_nxt_5_4_port, A2 => n27001, ZN => N859)
                           ;
   U2965 : AND2_X1 port map( A1 => regs_nxt_5_5_port, A2 => n27001, ZN => N860)
                           ;
   U2966 : AND2_X1 port map( A1 => regs_nxt_5_6_port, A2 => n27001, ZN => N861)
                           ;
   U2967 : AND2_X1 port map( A1 => regs_nxt_5_7_port, A2 => n27001, ZN => N862)
                           ;
   U2968 : AND2_X1 port map( A1 => regs_nxt_5_8_port, A2 => n27001, ZN => N863)
                           ;
   U2969 : AND2_X1 port map( A1 => regs_nxt_5_9_port, A2 => n27001, ZN => N864)
                           ;
   U2970 : AND2_X1 port map( A1 => regs_nxt_5_10_port, A2 => n27001, ZN => N865
                           );
   U2971 : AND2_X1 port map( A1 => regs_nxt_5_11_port, A2 => n27001, ZN => N866
                           );
   U2972 : AND2_X1 port map( A1 => regs_nxt_5_12_port, A2 => n27001, ZN => N867
                           );
   U2973 : AND2_X1 port map( A1 => regs_nxt_5_13_port, A2 => n27001, ZN => N868
                           );
   U2974 : AND2_X1 port map( A1 => regs_nxt_5_14_port, A2 => n27001, ZN => N869
                           );
   U2975 : AND2_X1 port map( A1 => regs_nxt_5_15_port, A2 => n27001, ZN => N870
                           );
   U2976 : AND2_X1 port map( A1 => regs_nxt_5_16_port, A2 => n27002, ZN => N871
                           );
   U2977 : AND2_X1 port map( A1 => regs_nxt_5_17_port, A2 => n27002, ZN => N872
                           );
   U2978 : AND2_X1 port map( A1 => regs_nxt_5_18_port, A2 => n27002, ZN => N873
                           );
   U2979 : AND2_X1 port map( A1 => regs_nxt_5_19_port, A2 => n27002, ZN => N874
                           );
   U2980 : AND2_X1 port map( A1 => regs_nxt_5_20_port, A2 => n27002, ZN => N875
                           );
   U2981 : AND2_X1 port map( A1 => regs_nxt_5_21_port, A2 => n27002, ZN => N876
                           );
   U2982 : AND2_X1 port map( A1 => regs_nxt_5_22_port, A2 => n27002, ZN => N877
                           );
   U2983 : AND2_X1 port map( A1 => regs_nxt_5_23_port, A2 => n27002, ZN => N878
                           );
   U2984 : AND2_X1 port map( A1 => regs_nxt_5_24_port, A2 => n27002, ZN => N879
                           );
   U2985 : AND2_X1 port map( A1 => regs_nxt_5_25_port, A2 => n27002, ZN => N880
                           );
   U2986 : AND2_X1 port map( A1 => regs_nxt_5_26_port, A2 => n27002, ZN => N881
                           );
   U2987 : AND2_X1 port map( A1 => regs_nxt_5_27_port, A2 => n27002, ZN => N882
                           );
   U2988 : AND2_X1 port map( A1 => regs_nxt_5_28_port, A2 => n27002, ZN => N883
                           );
   U2989 : AND2_X1 port map( A1 => regs_nxt_5_29_port, A2 => n27002, ZN => N884
                           );
   U2990 : AND2_X1 port map( A1 => regs_nxt_5_30_port, A2 => n27002, ZN => N885
                           );
   U2991 : AND2_X1 port map( A1 => regs_nxt_5_31_port, A2 => n27002, ZN => N886
                           );
   U2992 : AND2_X1 port map( A1 => regs_nxt_4_0_port, A2 => n27002, ZN => N887)
                           ;
   U2993 : AND2_X1 port map( A1 => regs_nxt_4_1_port, A2 => n27003, ZN => N888)
                           ;
   U2994 : AND2_X1 port map( A1 => regs_nxt_4_2_port, A2 => n27003, ZN => N889)
                           ;
   U2995 : AND2_X1 port map( A1 => regs_nxt_4_3_port, A2 => n27003, ZN => N890)
                           ;
   U2996 : AND2_X1 port map( A1 => regs_nxt_4_4_port, A2 => n27003, ZN => N891)
                           ;
   U2997 : AND2_X1 port map( A1 => regs_nxt_4_5_port, A2 => n27003, ZN => N892)
                           ;
   U2998 : AND2_X1 port map( A1 => regs_nxt_4_6_port, A2 => n27003, ZN => N893)
                           ;
   U2999 : AND2_X1 port map( A1 => regs_nxt_4_7_port, A2 => n27003, ZN => N894)
                           ;
   U3000 : AND2_X1 port map( A1 => regs_nxt_4_8_port, A2 => n27003, ZN => N895)
                           ;
   U3001 : AND2_X1 port map( A1 => regs_nxt_4_9_port, A2 => n27003, ZN => N896)
                           ;
   U3002 : AND2_X1 port map( A1 => regs_nxt_4_10_port, A2 => n27003, ZN => N897
                           );
   U3003 : AND2_X1 port map( A1 => regs_nxt_4_11_port, A2 => n27003, ZN => N898
                           );
   U3004 : AND2_X1 port map( A1 => regs_nxt_4_12_port, A2 => n27003, ZN => N899
                           );
   U3005 : AND2_X1 port map( A1 => regs_nxt_4_13_port, A2 => n27003, ZN => N900
                           );
   U3006 : AND2_X1 port map( A1 => regs_nxt_4_14_port, A2 => n27003, ZN => N901
                           );
   U3007 : AND2_X1 port map( A1 => regs_nxt_4_15_port, A2 => n27003, ZN => N902
                           );
   U3008 : AND2_X1 port map( A1 => regs_nxt_4_16_port, A2 => n27003, ZN => N903
                           );
   U3009 : AND2_X1 port map( A1 => regs_nxt_4_17_port, A2 => n27004, ZN => N904
                           );
   U3010 : AND2_X1 port map( A1 => regs_nxt_4_18_port, A2 => n27004, ZN => N905
                           );
   U3011 : AND2_X1 port map( A1 => regs_nxt_4_19_port, A2 => n27004, ZN => N906
                           );
   U3012 : AND2_X1 port map( A1 => regs_nxt_4_20_port, A2 => n27004, ZN => N907
                           );
   U3013 : AND2_X1 port map( A1 => regs_nxt_4_21_port, A2 => n26993, ZN => N908
                           );
   U3014 : AND2_X1 port map( A1 => regs_nxt_4_22_port, A2 => n26989, ZN => N909
                           );
   U3015 : AND2_X1 port map( A1 => regs_nxt_4_23_port, A2 => n26989, ZN => N910
                           );
   U3016 : AND2_X1 port map( A1 => regs_nxt_4_24_port, A2 => n26989, ZN => N911
                           );
   U3017 : AND2_X1 port map( A1 => regs_nxt_4_25_port, A2 => n26989, ZN => N912
                           );
   U3018 : AND2_X1 port map( A1 => regs_nxt_4_26_port, A2 => n26989, ZN => N913
                           );
   U3019 : AND2_X1 port map( A1 => regs_nxt_4_27_port, A2 => n26989, ZN => N914
                           );
   U3020 : AND2_X1 port map( A1 => regs_nxt_4_28_port, A2 => n26989, ZN => N915
                           );
   U3021 : AND2_X1 port map( A1 => regs_nxt_4_29_port, A2 => n26990, ZN => N916
                           );
   U3022 : AND2_X1 port map( A1 => regs_nxt_4_30_port, A2 => n26990, ZN => N917
                           );
   U3023 : AND2_X1 port map( A1 => regs_nxt_4_31_port, A2 => n26990, ZN => N918
                           );
   U3024 : AND2_X1 port map( A1 => regs_nxt_3_0_port, A2 => n26990, ZN => N919)
                           ;
   U3025 : AND2_X1 port map( A1 => regs_nxt_3_1_port, A2 => n26990, ZN => N920)
                           ;
   U3026 : AND2_X1 port map( A1 => regs_nxt_3_2_port, A2 => n26990, ZN => N921)
                           ;
   U3027 : AND2_X1 port map( A1 => regs_nxt_3_3_port, A2 => n26990, ZN => N922)
                           ;
   U3028 : AND2_X1 port map( A1 => regs_nxt_3_4_port, A2 => n26990, ZN => N923)
                           ;
   U3041 : AND2_X1 port map( A1 => regs_nxt_3_5_port, A2 => n26990, ZN => N924)
                           ;
   U3042 : AND2_X1 port map( A1 => regs_nxt_3_6_port, A2 => n26990, ZN => N925)
                           ;
   U3043 : AND2_X1 port map( A1 => regs_nxt_3_7_port, A2 => n26990, ZN => N926)
                           ;
   U3044 : AND2_X1 port map( A1 => regs_nxt_3_8_port, A2 => n26990, ZN => N927)
                           ;
   U3045 : AND2_X1 port map( A1 => regs_nxt_3_9_port, A2 => n26990, ZN => N928)
                           ;
   U3046 : AND2_X1 port map( A1 => regs_nxt_3_10_port, A2 => n26990, ZN => N929
                           );
   U3047 : AND2_X1 port map( A1 => regs_nxt_3_11_port, A2 => n26990, ZN => N930
                           );
   U3048 : AND2_X1 port map( A1 => regs_nxt_3_12_port, A2 => n26990, ZN => N931
                           );
   U3049 : AND2_X1 port map( A1 => regs_nxt_3_13_port, A2 => n26991, ZN => N932
                           );
   U3050 : AND2_X1 port map( A1 => regs_nxt_3_14_port, A2 => n26991, ZN => N933
                           );
   U3051 : AND2_X1 port map( A1 => regs_nxt_3_15_port, A2 => n26991, ZN => N934
                           );
   U3052 : AND2_X1 port map( A1 => regs_nxt_3_16_port, A2 => n26991, ZN => N935
                           );
   U3053 : AND2_X1 port map( A1 => regs_nxt_3_17_port, A2 => n26991, ZN => N936
                           );
   U3054 : AND2_X1 port map( A1 => regs_nxt_3_18_port, A2 => n26991, ZN => N937
                           );
   U3055 : AND2_X1 port map( A1 => regs_nxt_3_19_port, A2 => n26991, ZN => N938
                           );
   U3056 : AND2_X1 port map( A1 => regs_nxt_3_20_port, A2 => n26991, ZN => N939
                           );
   U3057 : AND2_X1 port map( A1 => regs_nxt_3_21_port, A2 => n26991, ZN => N940
                           );
   U3058 : AND2_X1 port map( A1 => regs_nxt_3_22_port, A2 => n26991, ZN => N941
                           );
   U3059 : AND2_X1 port map( A1 => regs_nxt_3_23_port, A2 => n26991, ZN => N942
                           );
   U3060 : AND2_X1 port map( A1 => regs_nxt_3_24_port, A2 => n26991, ZN => N943
                           );
   U3061 : AND2_X1 port map( A1 => regs_nxt_3_25_port, A2 => n26991, ZN => N944
                           );
   U3062 : AND2_X1 port map( A1 => regs_nxt_3_26_port, A2 => n26991, ZN => N945
                           );
   U3063 : AND2_X1 port map( A1 => regs_nxt_3_27_port, A2 => n26991, ZN => N946
                           );
   U3064 : AND2_X1 port map( A1 => regs_nxt_3_28_port, A2 => n26991, ZN => N947
                           );
   U3065 : AND2_X1 port map( A1 => regs_nxt_3_29_port, A2 => n26991, ZN => N948
                           );
   U3066 : AND2_X1 port map( A1 => regs_nxt_3_30_port, A2 => n26992, ZN => N949
                           );
   U3067 : AND2_X1 port map( A1 => regs_nxt_3_31_port, A2 => n26992, ZN => N950
                           );
   U3068 : AND2_X1 port map( A1 => regs_nxt_2_0_port, A2 => n26992, ZN => N951)
                           ;
   U3069 : AND2_X1 port map( A1 => regs_nxt_2_1_port, A2 => n26992, ZN => N952)
                           ;
   U3070 : AND2_X1 port map( A1 => regs_nxt_2_2_port, A2 => n26992, ZN => N953)
                           ;
   U3071 : AND2_X1 port map( A1 => regs_nxt_2_3_port, A2 => n26992, ZN => N954)
                           ;
   U3072 : AND2_X1 port map( A1 => regs_nxt_2_4_port, A2 => n26992, ZN => N955)
                           ;
   U3073 : AND2_X1 port map( A1 => regs_nxt_2_5_port, A2 => n26992, ZN => N956)
                           ;
   U3074 : AND2_X1 port map( A1 => regs_nxt_2_6_port, A2 => n26992, ZN => N957)
                           ;
   U3075 : AND2_X1 port map( A1 => regs_nxt_2_7_port, A2 => n26992, ZN => N958)
                           ;
   U3076 : AND2_X1 port map( A1 => regs_nxt_2_8_port, A2 => n26992, ZN => N959)
                           ;
   U3077 : AND2_X1 port map( A1 => regs_nxt_2_9_port, A2 => n26992, ZN => N960)
                           ;
   U3078 : AND2_X1 port map( A1 => regs_nxt_2_10_port, A2 => n26992, ZN => N961
                           );
   U3079 : AND2_X1 port map( A1 => regs_nxt_2_11_port, A2 => n26992, ZN => N962
                           );
   U3080 : AND2_X1 port map( A1 => regs_nxt_2_12_port, A2 => n26992, ZN => N963
                           );
   U3081 : AND2_X1 port map( A1 => regs_nxt_2_13_port, A2 => n26992, ZN => N964
                           );
   U3082 : AND2_X1 port map( A1 => regs_nxt_2_14_port, A2 => n26993, ZN => N965
                           );
   U3083 : AND2_X1 port map( A1 => regs_nxt_2_15_port, A2 => n26993, ZN => N966
                           );
   U3084 : AND2_X1 port map( A1 => regs_nxt_2_16_port, A2 => n26993, ZN => N967
                           );
   U3085 : AND2_X1 port map( A1 => regs_nxt_2_17_port, A2 => n26993, ZN => N968
                           );
   U3086 : AND2_X1 port map( A1 => regs_nxt_2_18_port, A2 => n26993, ZN => N969
                           );
   U3087 : AND2_X1 port map( A1 => regs_nxt_2_19_port, A2 => n26993, ZN => N970
                           );
   U3088 : AND2_X1 port map( A1 => regs_nxt_2_20_port, A2 => n26993, ZN => N971
                           );
   U3089 : AND2_X1 port map( A1 => regs_nxt_2_21_port, A2 => n26993, ZN => N972
                           );
   U3090 : AND2_X1 port map( A1 => regs_nxt_2_22_port, A2 => n26993, ZN => N973
                           );
   U3091 : AND2_X1 port map( A1 => regs_nxt_2_23_port, A2 => n26993, ZN => N974
                           );
   U3092 : AND2_X1 port map( A1 => regs_nxt_2_24_port, A2 => n26993, ZN => N975
                           );
   U3093 : AND2_X1 port map( A1 => regs_nxt_2_25_port, A2 => n26993, ZN => N976
                           );
   U3094 : AND2_X1 port map( A1 => regs_nxt_2_26_port, A2 => n26993, ZN => N977
                           );
   U3095 : AND2_X1 port map( A1 => regs_nxt_2_27_port, A2 => n26993, ZN => N978
                           );
   U3096 : AND2_X1 port map( A1 => regs_nxt_2_28_port, A2 => n26993, ZN => N979
                           );
   U3097 : AND2_X1 port map( A1 => regs_nxt_2_29_port, A2 => n26994, ZN => N980
                           );
   U3098 : AND2_X1 port map( A1 => regs_nxt_2_30_port, A2 => n26994, ZN => N981
                           );
   U3099 : AND2_X1 port map( A1 => regs_nxt_2_31_port, A2 => n26994, ZN => N982
                           );
   U3100 : AND2_X1 port map( A1 => regs_nxt_1_0_port, A2 => n26994, ZN => N983)
                           ;
   U3101 : AND2_X1 port map( A1 => regs_nxt_1_1_port, A2 => n26994, ZN => N984)
                           ;
   U3102 : AND2_X1 port map( A1 => regs_nxt_1_2_port, A2 => n26994, ZN => N985)
                           ;
   U3103 : AND2_X1 port map( A1 => regs_nxt_1_3_port, A2 => n26994, ZN => N986)
                           ;
   U3104 : AND2_X1 port map( A1 => regs_nxt_1_4_port, A2 => n26994, ZN => N987)
                           ;
   U3105 : AND2_X1 port map( A1 => regs_nxt_1_5_port, A2 => n26994, ZN => N988)
                           ;
   U3106 : AND2_X1 port map( A1 => regs_nxt_1_6_port, A2 => n26994, ZN => N989)
                           ;
   U3107 : AND2_X1 port map( A1 => regs_nxt_1_7_port, A2 => n26994, ZN => N990)
                           ;
   U3108 : AND2_X1 port map( A1 => regs_nxt_1_8_port, A2 => n26994, ZN => N991)
                           ;
   U3109 : AND2_X1 port map( A1 => regs_nxt_1_9_port, A2 => n26994, ZN => N992)
                           ;
   U3110 : AND2_X1 port map( A1 => regs_nxt_1_10_port, A2 => n26994, ZN => N993
                           );
   U3111 : AND2_X1 port map( A1 => regs_nxt_1_11_port, A2 => n26994, ZN => N994
                           );
   U3112 : AND2_X1 port map( A1 => regs_nxt_1_12_port, A2 => n26994, ZN => N995
                           );
   U3113 : AND2_X1 port map( A1 => regs_nxt_1_13_port, A2 => n26994, ZN => N996
                           );
   U3114 : AND2_X1 port map( A1 => regs_nxt_1_14_port, A2 => n26995, ZN => N997
                           );
   U3115 : AND2_X1 port map( A1 => regs_nxt_1_15_port, A2 => n26995, ZN => N998
                           );
   U3116 : AND2_X1 port map( A1 => regs_nxt_1_16_port, A2 => n26995, ZN => N999
                           );
   U3117 : AND2_X1 port map( A1 => regs_nxt_1_17_port, A2 => n27018, ZN => 
                           N1000);
   U3118 : AND2_X1 port map( A1 => regs_nxt_1_18_port, A2 => n27015, ZN => 
                           N1001);
   U3119 : AND2_X1 port map( A1 => regs_nxt_1_19_port, A2 => n27011, ZN => 
                           N1002);
   U3120 : AND2_X1 port map( A1 => regs_nxt_1_20_port, A2 => n27011, ZN => 
                           N1003);
   U3121 : AND2_X1 port map( A1 => regs_nxt_1_21_port, A2 => n27011, ZN => 
                           N1004);
   U3122 : AND2_X1 port map( A1 => regs_nxt_1_22_port, A2 => n27011, ZN => 
                           N1005);
   U3123 : AND2_X1 port map( A1 => regs_nxt_1_23_port, A2 => n27011, ZN => 
                           N1006);
   U3124 : AND2_X1 port map( A1 => regs_nxt_1_24_port, A2 => n27011, ZN => 
                           N1007);
   U3125 : AND2_X1 port map( A1 => regs_nxt_1_25_port, A2 => n27011, ZN => 
                           N1008);
   U3126 : AND2_X1 port map( A1 => regs_nxt_1_26_port, A2 => n27012, ZN => 
                           N1009);
   U3127 : AND2_X1 port map( A1 => regs_nxt_1_27_port, A2 => n27012, ZN => 
                           N1010);
   U3128 : AND2_X1 port map( A1 => regs_nxt_1_28_port, A2 => n27012, ZN => 
                           N1011);
   U3129 : AND2_X1 port map( A1 => regs_nxt_1_29_port, A2 => n27012, ZN => 
                           N1012);
   U3130 : AND2_X1 port map( A1 => regs_nxt_1_30_port, A2 => n27012, ZN => 
                           N1013);
   U3131 : AND2_X1 port map( A1 => regs_nxt_1_31_port, A2 => n27012, ZN => 
                           N1014);
   U3132 : AND2_X1 port map( A1 => regs_nxt_0_0_port, A2 => n27012, ZN => N1015
                           );
   U3133 : AND2_X1 port map( A1 => regs_nxt_0_1_port, A2 => n27012, ZN => N1016
                           );
   U3134 : AND2_X1 port map( A1 => regs_nxt_0_2_port, A2 => n27012, ZN => N1017
                           );
   U3135 : AND2_X1 port map( A1 => regs_nxt_0_3_port, A2 => n27012, ZN => N1018
                           );
   U3136 : AND2_X1 port map( A1 => regs_nxt_0_4_port, A2 => n27012, ZN => N1019
                           );
   U3137 : AND2_X1 port map( A1 => regs_nxt_0_5_port, A2 => n27012, ZN => N1020
                           );
   U3138 : AND2_X1 port map( A1 => regs_nxt_0_6_port, A2 => n27012, ZN => N1021
                           );
   U3139 : AND2_X1 port map( A1 => regs_nxt_0_7_port, A2 => n27012, ZN => N1022
                           );
   U3140 : AND2_X1 port map( A1 => regs_nxt_0_8_port, A2 => n27012, ZN => N1023
                           );
   U3141 : AND2_X1 port map( A1 => regs_nxt_0_9_port, A2 => n27012, ZN => N1024
                           );
   U3142 : AND2_X1 port map( A1 => regs_nxt_0_10_port, A2 => n27013, ZN => 
                           N1025);
   U3143 : AND2_X1 port map( A1 => regs_nxt_0_11_port, A2 => n27013, ZN => 
                           N1026);
   U3144 : AND2_X1 port map( A1 => regs_nxt_0_12_port, A2 => n27013, ZN => 
                           N1027);
   U3145 : AND2_X1 port map( A1 => regs_nxt_0_13_port, A2 => n27013, ZN => 
                           N1028);
   U3146 : AND2_X1 port map( A1 => regs_nxt_0_14_port, A2 => n27013, ZN => 
                           N1029);
   U3147 : AND2_X1 port map( A1 => regs_nxt_0_15_port, A2 => n27013, ZN => 
                           N1030);
   U3148 : AND2_X1 port map( A1 => regs_nxt_0_16_port, A2 => n27013, ZN => 
                           N1031);
   U3149 : AND2_X1 port map( A1 => regs_nxt_0_17_port, A2 => n27013, ZN => 
                           N1032);
   U3150 : AND2_X1 port map( A1 => regs_nxt_0_18_port, A2 => n27013, ZN => 
                           N1033);
   U3151 : AND2_X1 port map( A1 => regs_nxt_0_19_port, A2 => n27013, ZN => 
                           N1034);
   U3152 : AND2_X1 port map( A1 => regs_nxt_0_20_port, A2 => n27013, ZN => 
                           N1035);
   U3153 : AND2_X1 port map( A1 => regs_nxt_0_21_port, A2 => n27013, ZN => 
                           N1036);
   U3154 : AND2_X1 port map( A1 => regs_nxt_0_22_port, A2 => n27013, ZN => 
                           N1037);
   U3155 : AND2_X1 port map( A1 => regs_nxt_0_23_port, A2 => n27013, ZN => 
                           N1038);
   U3156 : AND2_X1 port map( A1 => regs_nxt_0_24_port, A2 => n27013, ZN => 
                           N1039);
   U3157 : AND2_X1 port map( A1 => regs_nxt_0_25_port, A2 => n27013, ZN => 
                           N1040);
   U3158 : AND2_X1 port map( A1 => regs_nxt_0_26_port, A2 => n27014, ZN => 
                           N1041);
   U3159 : AND2_X1 port map( A1 => regs_nxt_0_27_port, A2 => n27014, ZN => 
                           N1042);
   U3160 : AND2_X1 port map( A1 => regs_nxt_0_28_port, A2 => n27014, ZN => 
                           N1043);
   U3161 : AND2_X1 port map( A1 => regs_nxt_0_29_port, A2 => n27014, ZN => 
                           N1044);
   U3162 : AND2_X1 port map( A1 => regs_nxt_0_30_port, A2 => n27014, ZN => 
                           N1045);
   U3163 : AND2_X1 port map( A1 => regs_nxt_0_31_port, A2 => n27014, ZN => 
                           N1046);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity add4_NBIT32 is

   port( A : in std_logic_vector (31 downto 0);  res : out std_logic_vector (31
         downto 0));

end add4_NBIT32;

architecture SYN_beh of add4_NBIT32 is

   component add4_NBIT32_DW01_add_0_DW01_add_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1627 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   add_17 : add4_NBIT32_DW01_add_0_DW01_add_2 port map( A(31) => A(31), A(30) 
                           => A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => n3, B(30) => n3, 
                           B(29) => n3, B(28) => n3, B(27) => n3, B(26) => n3, 
                           B(25) => n3, B(24) => n3, B(23) => n3, B(22) => n3, 
                           B(21) => n3, B(20) => n3, B(19) => n3, B(18) => n3, 
                           B(17) => n3, B(16) => n3, B(15) => n3, B(14) => n3, 
                           B(13) => n3, B(12) => n3, B(11) => n3, B(10) => n3, 
                           B(9) => n3, B(8) => n3, B(7) => n3, B(6) => n3, B(5)
                           => n3, B(4) => n3, B(3) => n3, B(2) => n2, B(1) => 
                           n1, B(0) => n1, CI => n3, SUM(31) => res(31), 
                           SUM(30) => res(30), SUM(29) => res(29), SUM(28) => 
                           res(28), SUM(27) => res(27), SUM(26) => res(26), 
                           SUM(25) => res(25), SUM(24) => res(24), SUM(23) => 
                           res(23), SUM(22) => res(22), SUM(21) => res(21), 
                           SUM(20) => res(20), SUM(19) => res(19), SUM(18) => 
                           res(18), SUM(17) => res(17), SUM(16) => res(16), 
                           SUM(15) => res(15), SUM(14) => res(14), SUM(13) => 
                           res(13), SUM(12) => res(12), SUM(11) => res(11), 
                           SUM(10) => res(10), SUM(9) => res(9), SUM(8) => 
                           res(8), SUM(7) => res(7), SUM(6) => res(6), SUM(5) 
                           => res(5), SUM(4) => res(4), SUM(3) => res(3), 
                           SUM(2) => res(2), SUM(1) => res(1), SUM(0) => res(0)
                           , CO => n_1627);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity WBU_N32 is

   port( ALU_OUT, LOAD, NPC_REG_in, RT_REG_in : in std_logic_vector (31 downto 
         0);  IS_JAL, ALUOUT_OR_LOAD : in std_logic;  RF_ADDR, RF_DATA : out 
         std_logic_vector (31 downto 0));

end WBU_N32;

architecture SYN_STRUCTURAL of WBU_N32 is

   component mux21_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   signal alu_lmd_s_9_port, alu_lmd_s_8_port, alu_lmd_s_7_port, 
      alu_lmd_s_6_port, alu_lmd_s_5_port, alu_lmd_s_4_port, alu_lmd_s_3_port, 
      alu_lmd_s_31_port, alu_lmd_s_30_port, alu_lmd_s_2_port, alu_lmd_s_29_port
      , alu_lmd_s_28_port, alu_lmd_s_27_port, alu_lmd_s_26_port, 
      alu_lmd_s_25_port, alu_lmd_s_24_port, alu_lmd_s_23_port, 
      alu_lmd_s_22_port, alu_lmd_s_21_port, alu_lmd_s_20_port, alu_lmd_s_1_port
      , alu_lmd_s_19_port, alu_lmd_s_18_port, alu_lmd_s_17_port, 
      alu_lmd_s_16_port, alu_lmd_s_15_port, alu_lmd_s_14_port, 
      alu_lmd_s_13_port, alu_lmd_s_12_port, alu_lmd_s_11_port, 
      alu_lmd_s_10_port, alu_lmd_s_0_port, n33, n34 : std_logic;

begin
   
   alu_lmd_mux : mux21_NBIT32_3 port map( A(31) => ALU_OUT(31), A(30) => 
                           ALU_OUT(30), A(29) => ALU_OUT(29), A(28) => 
                           ALU_OUT(28), A(27) => ALU_OUT(27), A(26) => 
                           ALU_OUT(26), A(25) => ALU_OUT(25), A(24) => 
                           ALU_OUT(24), A(23) => ALU_OUT(23), A(22) => 
                           ALU_OUT(22), A(21) => ALU_OUT(21), A(20) => 
                           ALU_OUT(20), A(19) => ALU_OUT(19), A(18) => 
                           ALU_OUT(18), A(17) => ALU_OUT(17), A(16) => 
                           ALU_OUT(16), A(15) => ALU_OUT(15), A(14) => 
                           ALU_OUT(14), A(13) => ALU_OUT(13), A(12) => 
                           ALU_OUT(12), A(11) => ALU_OUT(11), A(10) => 
                           ALU_OUT(10), A(9) => ALU_OUT(9), A(8) => ALU_OUT(8),
                           A(7) => ALU_OUT(7), A(6) => ALU_OUT(6), A(5) => 
                           ALU_OUT(5), A(4) => ALU_OUT(4), A(3) => ALU_OUT(3), 
                           A(2) => ALU_OUT(2), A(1) => ALU_OUT(1), A(0) => 
                           ALU_OUT(0), B(31) => LOAD(31), B(30) => LOAD(30), 
                           B(29) => LOAD(29), B(28) => LOAD(28), B(27) => 
                           LOAD(27), B(26) => LOAD(26), B(25) => LOAD(25), 
                           B(24) => LOAD(24), B(23) => LOAD(23), B(22) => 
                           LOAD(22), B(21) => LOAD(21), B(20) => LOAD(20), 
                           B(19) => LOAD(19), B(18) => LOAD(18), B(17) => 
                           LOAD(17), B(16) => LOAD(16), B(15) => LOAD(15), 
                           B(14) => LOAD(14), B(13) => LOAD(13), B(12) => 
                           LOAD(12), B(11) => LOAD(11), B(10) => LOAD(10), B(9)
                           => LOAD(9), B(8) => LOAD(8), B(7) => LOAD(7), B(6) 
                           => LOAD(6), B(5) => LOAD(5), B(4) => LOAD(4), B(3) 
                           => LOAD(3), B(2) => LOAD(2), B(1) => LOAD(1), B(0) 
                           => LOAD(0), sel => ALUOUT_OR_LOAD, muxout(31) => 
                           alu_lmd_s_31_port, muxout(30) => alu_lmd_s_30_port, 
                           muxout(29) => alu_lmd_s_29_port, muxout(28) => 
                           alu_lmd_s_28_port, muxout(27) => alu_lmd_s_27_port, 
                           muxout(26) => alu_lmd_s_26_port, muxout(25) => 
                           alu_lmd_s_25_port, muxout(24) => alu_lmd_s_24_port, 
                           muxout(23) => alu_lmd_s_23_port, muxout(22) => 
                           alu_lmd_s_22_port, muxout(21) => alu_lmd_s_21_port, 
                           muxout(20) => alu_lmd_s_20_port, muxout(19) => 
                           alu_lmd_s_19_port, muxout(18) => alu_lmd_s_18_port, 
                           muxout(17) => alu_lmd_s_17_port, muxout(16) => 
                           alu_lmd_s_16_port, muxout(15) => alu_lmd_s_15_port, 
                           muxout(14) => alu_lmd_s_14_port, muxout(13) => 
                           alu_lmd_s_13_port, muxout(12) => alu_lmd_s_12_port, 
                           muxout(11) => alu_lmd_s_11_port, muxout(10) => 
                           alu_lmd_s_10_port, muxout(9) => alu_lmd_s_9_port, 
                           muxout(8) => alu_lmd_s_8_port, muxout(7) => 
                           alu_lmd_s_7_port, muxout(6) => alu_lmd_s_6_port, 
                           muxout(5) => alu_lmd_s_5_port, muxout(4) => 
                           alu_lmd_s_4_port, muxout(3) => alu_lmd_s_3_port, 
                           muxout(2) => alu_lmd_s_2_port, muxout(1) => 
                           alu_lmd_s_1_port, muxout(0) => alu_lmd_s_0_port);
   addr_mux : mux21_NBIT32_2 port map( A(31) => n34, A(30) => n34, A(29) => n34
                           , A(28) => n34, A(27) => n34, A(26) => n34, A(25) =>
                           n34, A(24) => n34, A(23) => n34, A(22) => n34, A(21)
                           => n34, A(20) => n34, A(19) => n34, A(18) => n34, 
                           A(17) => n34, A(16) => n34, A(15) => n34, A(14) => 
                           n34, A(13) => n34, A(12) => n34, A(11) => n34, A(10)
                           => n34, A(9) => n34, A(8) => n34, A(7) => n34, A(6) 
                           => n34, A(5) => n34, A(4) => n33, A(3) => n33, A(2) 
                           => n33, A(1) => n33, A(0) => n33, B(31) => 
                           RT_REG_in(31), B(30) => RT_REG_in(30), B(29) => 
                           RT_REG_in(29), B(28) => RT_REG_in(28), B(27) => 
                           RT_REG_in(27), B(26) => RT_REG_in(26), B(25) => 
                           RT_REG_in(25), B(24) => RT_REG_in(24), B(23) => 
                           RT_REG_in(23), B(22) => RT_REG_in(22), B(21) => 
                           RT_REG_in(21), B(20) => RT_REG_in(20), B(19) => 
                           RT_REG_in(19), B(18) => RT_REG_in(18), B(17) => 
                           RT_REG_in(17), B(16) => RT_REG_in(16), B(15) => 
                           RT_REG_in(15), B(14) => RT_REG_in(14), B(13) => 
                           RT_REG_in(13), B(12) => RT_REG_in(12), B(11) => 
                           RT_REG_in(11), B(10) => RT_REG_in(10), B(9) => 
                           RT_REG_in(9), B(8) => RT_REG_in(8), B(7) => 
                           RT_REG_in(7), B(6) => RT_REG_in(6), B(5) => 
                           RT_REG_in(5), B(4) => RT_REG_in(4), B(3) => 
                           RT_REG_in(3), B(2) => RT_REG_in(2), B(1) => 
                           RT_REG_in(1), B(0) => RT_REG_in(0), sel => IS_JAL, 
                           muxout(31) => RF_ADDR(31), muxout(30) => RF_ADDR(30)
                           , muxout(29) => RF_ADDR(29), muxout(28) => 
                           RF_ADDR(28), muxout(27) => RF_ADDR(27), muxout(26) 
                           => RF_ADDR(26), muxout(25) => RF_ADDR(25), 
                           muxout(24) => RF_ADDR(24), muxout(23) => RF_ADDR(23)
                           , muxout(22) => RF_ADDR(22), muxout(21) => 
                           RF_ADDR(21), muxout(20) => RF_ADDR(20), muxout(19) 
                           => RF_ADDR(19), muxout(18) => RF_ADDR(18), 
                           muxout(17) => RF_ADDR(17), muxout(16) => RF_ADDR(16)
                           , muxout(15) => RF_ADDR(15), muxout(14) => 
                           RF_ADDR(14), muxout(13) => RF_ADDR(13), muxout(12) 
                           => RF_ADDR(12), muxout(11) => RF_ADDR(11), 
                           muxout(10) => RF_ADDR(10), muxout(9) => RF_ADDR(9), 
                           muxout(8) => RF_ADDR(8), muxout(7) => RF_ADDR(7), 
                           muxout(6) => RF_ADDR(6), muxout(5) => RF_ADDR(5), 
                           muxout(4) => RF_ADDR(4), muxout(3) => RF_ADDR(3), 
                           muxout(2) => RF_ADDR(2), muxout(1) => RF_ADDR(1), 
                           muxout(0) => RF_ADDR(0));
   data_mux : mux21_NBIT32_1 port map( A(31) => NPC_REG_in(31), A(30) => 
                           NPC_REG_in(30), A(29) => NPC_REG_in(29), A(28) => 
                           NPC_REG_in(28), A(27) => NPC_REG_in(27), A(26) => 
                           NPC_REG_in(26), A(25) => NPC_REG_in(25), A(24) => 
                           NPC_REG_in(24), A(23) => NPC_REG_in(23), A(22) => 
                           NPC_REG_in(22), A(21) => NPC_REG_in(21), A(20) => 
                           NPC_REG_in(20), A(19) => NPC_REG_in(19), A(18) => 
                           NPC_REG_in(18), A(17) => NPC_REG_in(17), A(16) => 
                           NPC_REG_in(16), A(15) => NPC_REG_in(15), A(14) => 
                           NPC_REG_in(14), A(13) => NPC_REG_in(13), A(12) => 
                           NPC_REG_in(12), A(11) => NPC_REG_in(11), A(10) => 
                           NPC_REG_in(10), A(9) => NPC_REG_in(9), A(8) => 
                           NPC_REG_in(8), A(7) => NPC_REG_in(7), A(6) => 
                           NPC_REG_in(6), A(5) => NPC_REG_in(5), A(4) => 
                           NPC_REG_in(4), A(3) => NPC_REG_in(3), A(2) => 
                           NPC_REG_in(2), A(1) => NPC_REG_in(1), A(0) => 
                           NPC_REG_in(0), B(31) => alu_lmd_s_31_port, B(30) => 
                           alu_lmd_s_30_port, B(29) => alu_lmd_s_29_port, B(28)
                           => alu_lmd_s_28_port, B(27) => alu_lmd_s_27_port, 
                           B(26) => alu_lmd_s_26_port, B(25) => 
                           alu_lmd_s_25_port, B(24) => alu_lmd_s_24_port, B(23)
                           => alu_lmd_s_23_port, B(22) => alu_lmd_s_22_port, 
                           B(21) => alu_lmd_s_21_port, B(20) => 
                           alu_lmd_s_20_port, B(19) => alu_lmd_s_19_port, B(18)
                           => alu_lmd_s_18_port, B(17) => alu_lmd_s_17_port, 
                           B(16) => alu_lmd_s_16_port, B(15) => 
                           alu_lmd_s_15_port, B(14) => alu_lmd_s_14_port, B(13)
                           => alu_lmd_s_13_port, B(12) => alu_lmd_s_12_port, 
                           B(11) => alu_lmd_s_11_port, B(10) => 
                           alu_lmd_s_10_port, B(9) => alu_lmd_s_9_port, B(8) =>
                           alu_lmd_s_8_port, B(7) => alu_lmd_s_7_port, B(6) => 
                           alu_lmd_s_6_port, B(5) => alu_lmd_s_5_port, B(4) => 
                           alu_lmd_s_4_port, B(3) => alu_lmd_s_3_port, B(2) => 
                           alu_lmd_s_2_port, B(1) => alu_lmd_s_1_port, B(0) => 
                           alu_lmd_s_0_port, sel => IS_JAL, muxout(31) => 
                           RF_DATA(31), muxout(30) => RF_DATA(30), muxout(29) 
                           => RF_DATA(29), muxout(28) => RF_DATA(28), 
                           muxout(27) => RF_DATA(27), muxout(26) => RF_DATA(26)
                           , muxout(25) => RF_DATA(25), muxout(24) => 
                           RF_DATA(24), muxout(23) => RF_DATA(23), muxout(22) 
                           => RF_DATA(22), muxout(21) => RF_DATA(21), 
                           muxout(20) => RF_DATA(20), muxout(19) => RF_DATA(19)
                           , muxout(18) => RF_DATA(18), muxout(17) => 
                           RF_DATA(17), muxout(16) => RF_DATA(16), muxout(15) 
                           => RF_DATA(15), muxout(14) => RF_DATA(14), 
                           muxout(13) => RF_DATA(13), muxout(12) => RF_DATA(12)
                           , muxout(11) => RF_DATA(11), muxout(10) => 
                           RF_DATA(10), muxout(9) => RF_DATA(9), muxout(8) => 
                           RF_DATA(8), muxout(7) => RF_DATA(7), muxout(6) => 
                           RF_DATA(6), muxout(5) => RF_DATA(5), muxout(4) => 
                           RF_DATA(4), muxout(3) => RF_DATA(3), muxout(2) => 
                           RF_DATA(2), muxout(1) => RF_DATA(1), muxout(0) => 
                           RF_DATA(0));
   n33 <= '1';
   n34 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MU_N32 is

   port( CLK, RST, LMD_EN : in std_logic;  ALU_RESULT, RT_REG_in, NPC_REG_in, 
         LMD_LATCH_in : in std_logic_vector (31 downto 0);  LMD_LATCH_out, 
         ALU_REG_out, RT_REG_out, NPC_REG_out : out std_logic_vector (31 downto
         0));

end MU_N32;

architecture SYN_structural of MU_N32 is

   component reg_N32_1
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_2
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_3
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_4
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   signal n15 : std_logic;

begin
   
   LMD_REG : reg_N32_4 port map( clk => CLK, rst => RST, en => LMD_EN, A(31) =>
                           LMD_LATCH_in(31), A(30) => LMD_LATCH_in(30), A(29) 
                           => LMD_LATCH_in(29), A(28) => LMD_LATCH_in(28), 
                           A(27) => LMD_LATCH_in(27), A(26) => LMD_LATCH_in(26)
                           , A(25) => LMD_LATCH_in(25), A(24) => 
                           LMD_LATCH_in(24), A(23) => LMD_LATCH_in(23), A(22) 
                           => LMD_LATCH_in(22), A(21) => LMD_LATCH_in(21), 
                           A(20) => LMD_LATCH_in(20), A(19) => LMD_LATCH_in(19)
                           , A(18) => LMD_LATCH_in(18), A(17) => 
                           LMD_LATCH_in(17), A(16) => LMD_LATCH_in(16), A(15) 
                           => LMD_LATCH_in(15), A(14) => LMD_LATCH_in(14), 
                           A(13) => LMD_LATCH_in(13), A(12) => LMD_LATCH_in(12)
                           , A(11) => LMD_LATCH_in(11), A(10) => 
                           LMD_LATCH_in(10), A(9) => LMD_LATCH_in(9), A(8) => 
                           LMD_LATCH_in(8), A(7) => LMD_LATCH_in(7), A(6) => 
                           LMD_LATCH_in(6), A(5) => LMD_LATCH_in(5), A(4) => 
                           LMD_LATCH_in(4), A(3) => LMD_LATCH_in(3), A(2) => 
                           LMD_LATCH_in(2), A(1) => LMD_LATCH_in(1), A(0) => 
                           LMD_LATCH_in(0), Y(31) => LMD_LATCH_out(31), Y(30) 
                           => LMD_LATCH_out(30), Y(29) => LMD_LATCH_out(29), 
                           Y(28) => LMD_LATCH_out(28), Y(27) => 
                           LMD_LATCH_out(27), Y(26) => LMD_LATCH_out(26), Y(25)
                           => LMD_LATCH_out(25), Y(24) => LMD_LATCH_out(24), 
                           Y(23) => LMD_LATCH_out(23), Y(22) => 
                           LMD_LATCH_out(22), Y(21) => LMD_LATCH_out(21), Y(20)
                           => LMD_LATCH_out(20), Y(19) => LMD_LATCH_out(19), 
                           Y(18) => LMD_LATCH_out(18), Y(17) => 
                           LMD_LATCH_out(17), Y(16) => LMD_LATCH_out(16), Y(15)
                           => LMD_LATCH_out(15), Y(14) => LMD_LATCH_out(14), 
                           Y(13) => LMD_LATCH_out(13), Y(12) => 
                           LMD_LATCH_out(12), Y(11) => LMD_LATCH_out(11), Y(10)
                           => LMD_LATCH_out(10), Y(9) => LMD_LATCH_out(9), Y(8)
                           => LMD_LATCH_out(8), Y(7) => LMD_LATCH_out(7), Y(6) 
                           => LMD_LATCH_out(6), Y(5) => LMD_LATCH_out(5), Y(4) 
                           => LMD_LATCH_out(4), Y(3) => LMD_LATCH_out(3), Y(2) 
                           => LMD_LATCH_out(2), Y(1) => LMD_LATCH_out(1), Y(0) 
                           => LMD_LATCH_out(0));
   ALU_OUT_REG_1 : reg_N32_3 port map( clk => CLK, rst => RST, en => n15, A(31)
                           => ALU_RESULT(31), A(30) => ALU_RESULT(30), A(29) =>
                           ALU_RESULT(29), A(28) => ALU_RESULT(28), A(27) => 
                           ALU_RESULT(27), A(26) => ALU_RESULT(26), A(25) => 
                           ALU_RESULT(25), A(24) => ALU_RESULT(24), A(23) => 
                           ALU_RESULT(23), A(22) => ALU_RESULT(22), A(21) => 
                           ALU_RESULT(21), A(20) => ALU_RESULT(20), A(19) => 
                           ALU_RESULT(19), A(18) => ALU_RESULT(18), A(17) => 
                           ALU_RESULT(17), A(16) => ALU_RESULT(16), A(15) => 
                           ALU_RESULT(15), A(14) => ALU_RESULT(14), A(13) => 
                           ALU_RESULT(13), A(12) => ALU_RESULT(12), A(11) => 
                           ALU_RESULT(11), A(10) => ALU_RESULT(10), A(9) => 
                           ALU_RESULT(9), A(8) => ALU_RESULT(8), A(7) => 
                           ALU_RESULT(7), A(6) => ALU_RESULT(6), A(5) => 
                           ALU_RESULT(5), A(4) => ALU_RESULT(4), A(3) => 
                           ALU_RESULT(3), A(2) => ALU_RESULT(2), A(1) => 
                           ALU_RESULT(1), A(0) => ALU_RESULT(0), Y(31) => 
                           ALU_REG_out(31), Y(30) => ALU_REG_out(30), Y(29) => 
                           ALU_REG_out(29), Y(28) => ALU_REG_out(28), Y(27) => 
                           ALU_REG_out(27), Y(26) => ALU_REG_out(26), Y(25) => 
                           ALU_REG_out(25), Y(24) => ALU_REG_out(24), Y(23) => 
                           ALU_REG_out(23), Y(22) => ALU_REG_out(22), Y(21) => 
                           ALU_REG_out(21), Y(20) => ALU_REG_out(20), Y(19) => 
                           ALU_REG_out(19), Y(18) => ALU_REG_out(18), Y(17) => 
                           ALU_REG_out(17), Y(16) => ALU_REG_out(16), Y(15) => 
                           ALU_REG_out(15), Y(14) => ALU_REG_out(14), Y(13) => 
                           ALU_REG_out(13), Y(12) => ALU_REG_out(12), Y(11) => 
                           ALU_REG_out(11), Y(10) => ALU_REG_out(10), Y(9) => 
                           ALU_REG_out(9), Y(8) => ALU_REG_out(8), Y(7) => 
                           ALU_REG_out(7), Y(6) => ALU_REG_out(6), Y(5) => 
                           ALU_REG_out(5), Y(4) => ALU_REG_out(4), Y(3) => 
                           ALU_REG_out(3), Y(2) => ALU_REG_out(2), Y(1) => 
                           ALU_REG_out(1), Y(0) => ALU_REG_out(0));
   RT_REG_3 : reg_N32_2 port map( clk => CLK, rst => RST, en => n15, A(31) => 
                           RT_REG_in(31), A(30) => RT_REG_in(30), A(29) => 
                           RT_REG_in(29), A(28) => RT_REG_in(28), A(27) => 
                           RT_REG_in(27), A(26) => RT_REG_in(26), A(25) => 
                           RT_REG_in(25), A(24) => RT_REG_in(24), A(23) => 
                           RT_REG_in(23), A(22) => RT_REG_in(22), A(21) => 
                           RT_REG_in(21), A(20) => RT_REG_in(20), A(19) => 
                           RT_REG_in(19), A(18) => RT_REG_in(18), A(17) => 
                           RT_REG_in(17), A(16) => RT_REG_in(16), A(15) => 
                           RT_REG_in(15), A(14) => RT_REG_in(14), A(13) => 
                           RT_REG_in(13), A(12) => RT_REG_in(12), A(11) => 
                           RT_REG_in(11), A(10) => RT_REG_in(10), A(9) => 
                           RT_REG_in(9), A(8) => RT_REG_in(8), A(7) => 
                           RT_REG_in(7), A(6) => RT_REG_in(6), A(5) => 
                           RT_REG_in(5), A(4) => RT_REG_in(4), A(3) => 
                           RT_REG_in(3), A(2) => RT_REG_in(2), A(1) => 
                           RT_REG_in(1), A(0) => RT_REG_in(0), Y(31) => 
                           RT_REG_out(31), Y(30) => RT_REG_out(30), Y(29) => 
                           RT_REG_out(29), Y(28) => RT_REG_out(28), Y(27) => 
                           RT_REG_out(27), Y(26) => RT_REG_out(26), Y(25) => 
                           RT_REG_out(25), Y(24) => RT_REG_out(24), Y(23) => 
                           RT_REG_out(23), Y(22) => RT_REG_out(22), Y(21) => 
                           RT_REG_out(21), Y(20) => RT_REG_out(20), Y(19) => 
                           RT_REG_out(19), Y(18) => RT_REG_out(18), Y(17) => 
                           RT_REG_out(17), Y(16) => RT_REG_out(16), Y(15) => 
                           RT_REG_out(15), Y(14) => RT_REG_out(14), Y(13) => 
                           RT_REG_out(13), Y(12) => RT_REG_out(12), Y(11) => 
                           RT_REG_out(11), Y(10) => RT_REG_out(10), Y(9) => 
                           RT_REG_out(9), Y(8) => RT_REG_out(8), Y(7) => 
                           RT_REG_out(7), Y(6) => RT_REG_out(6), Y(5) => 
                           RT_REG_out(5), Y(4) => RT_REG_out(4), Y(3) => 
                           RT_REG_out(3), Y(2) => RT_REG_out(2), Y(1) => 
                           RT_REG_out(1), Y(0) => RT_REG_out(0));
   JAL_NPC_m : reg_N32_1 port map( clk => CLK, rst => RST, en => n15, A(31) => 
                           NPC_REG_in(31), A(30) => NPC_REG_in(30), A(29) => 
                           NPC_REG_in(29), A(28) => NPC_REG_in(28), A(27) => 
                           NPC_REG_in(27), A(26) => NPC_REG_in(26), A(25) => 
                           NPC_REG_in(25), A(24) => NPC_REG_in(24), A(23) => 
                           NPC_REG_in(23), A(22) => NPC_REG_in(22), A(21) => 
                           NPC_REG_in(21), A(20) => NPC_REG_in(20), A(19) => 
                           NPC_REG_in(19), A(18) => NPC_REG_in(18), A(17) => 
                           NPC_REG_in(17), A(16) => NPC_REG_in(16), A(15) => 
                           NPC_REG_in(15), A(14) => NPC_REG_in(14), A(13) => 
                           NPC_REG_in(13), A(12) => NPC_REG_in(12), A(11) => 
                           NPC_REG_in(11), A(10) => NPC_REG_in(10), A(9) => 
                           NPC_REG_in(9), A(8) => NPC_REG_in(8), A(7) => 
                           NPC_REG_in(7), A(6) => NPC_REG_in(6), A(5) => 
                           NPC_REG_in(5), A(4) => NPC_REG_in(4), A(3) => 
                           NPC_REG_in(3), A(2) => NPC_REG_in(2), A(1) => 
                           NPC_REG_in(1), A(0) => NPC_REG_in(0), Y(31) => 
                           NPC_REG_out(31), Y(30) => NPC_REG_out(30), Y(29) => 
                           NPC_REG_out(29), Y(28) => NPC_REG_out(28), Y(27) => 
                           NPC_REG_out(27), Y(26) => NPC_REG_out(26), Y(25) => 
                           NPC_REG_out(25), Y(24) => NPC_REG_out(24), Y(23) => 
                           NPC_REG_out(23), Y(22) => NPC_REG_out(22), Y(21) => 
                           NPC_REG_out(21), Y(20) => NPC_REG_out(20), Y(19) => 
                           NPC_REG_out(19), Y(18) => NPC_REG_out(18), Y(17) => 
                           NPC_REG_out(17), Y(16) => NPC_REG_out(16), Y(15) => 
                           NPC_REG_out(15), Y(14) => NPC_REG_out(14), Y(13) => 
                           NPC_REG_out(13), Y(12) => NPC_REG_out(12), Y(11) => 
                           NPC_REG_out(11), Y(10) => NPC_REG_out(10), Y(9) => 
                           NPC_REG_out(9), Y(8) => NPC_REG_out(8), Y(7) => 
                           NPC_REG_out(7), Y(6) => NPC_REG_out(6), Y(5) => 
                           NPC_REG_out(5), Y(4) => NPC_REG_out(4), Y(3) => 
                           NPC_REG_out(3), Y(2) => NPC_REG_out(2), Y(1) => 
                           NPC_REG_out(1), Y(0) => NPC_REG_out(0));
   n15 <= '1';

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity EXU_N32 is

   port( CLK, RST, MUXA_SEL, MUXB_SEL, ZERO_EN, ZERO_SEL, ALUOUT_EN, SHIFT2_EN 
         : in std_logic;  ALU_FUNC : in std_logic_vector (0 to 3);  NPC_REG, 
         A_REG, B_REG, RT_REG, IMM_REG, PC_4 : in std_logic_vector (31 downto 
         0);  ZERO : out std_logic;  BRANC_ADDR, ALU_OUT, RT_REG_OUT, NPC_OUT :
         out std_logic_vector (31 downto 0));

end EXU_N32;

architecture SYN_structural of EXU_N32 is

   component reg_N32_5
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_6
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_7
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component is_zero_NBIT32
      port( A : in std_logic_vector (31 downto 0);  BEQZ_OR_BNEZ, EN : in 
            std_logic;  res : out std_logic);
   end component;
   
   component ALU_N32
      port( FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux21_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   signal ZERO_port, op_1_s_31_port, op_1_s_30_port, op_1_s_29_port, 
      op_1_s_28_port, op_1_s_27_port, op_1_s_26_port, op_1_s_25_port, 
      op_1_s_24_port, op_1_s_23_port, op_1_s_22_port, op_1_s_21_port, 
      op_1_s_20_port, op_1_s_19_port, op_1_s_18_port, op_1_s_17_port, 
      op_1_s_16_port, op_1_s_15_port, op_1_s_14_port, op_1_s_13_port, 
      op_1_s_12_port, op_1_s_11_port, op_1_s_10_port, op_1_s_9_port, 
      op_1_s_8_port, op_1_s_7_port, op_1_s_6_port, op_1_s_5_port, op_1_s_4_port
      , op_1_s_3_port, op_1_s_2_port, op_1_s_1_port, op_1_s_0_port, 
      op_2_s_31_port, op_2_s_30_port, op_2_s_29_port, op_2_s_28_port, 
      op_2_s_27_port, op_2_s_26_port, op_2_s_25_port, op_2_s_24_port, 
      op_2_s_23_port, op_2_s_22_port, op_2_s_21_port, op_2_s_20_port, 
      op_2_s_19_port, op_2_s_18_port, op_2_s_17_port, op_2_s_16_port, 
      op_2_s_15_port, op_2_s_14_port, op_2_s_13_port, op_2_s_12_port, 
      op_2_s_11_port, op_2_s_10_port, op_2_s_9_port, op_2_s_8_port, 
      op_2_s_7_port, op_2_s_6_port, op_2_s_5_port, op_2_s_4_port, op_2_s_3_port
      , op_2_s_2_port, op_2_s_1_port, op_2_s_0_port, alu_out_s_31_port, 
      alu_out_s_30_port, alu_out_s_29_port, alu_out_s_28_port, 
      alu_out_s_27_port, alu_out_s_26_port, alu_out_s_25_port, 
      alu_out_s_24_port, alu_out_s_23_port, alu_out_s_22_port, 
      alu_out_s_21_port, alu_out_s_20_port, alu_out_s_19_port, 
      alu_out_s_18_port, alu_out_s_17_port, alu_out_s_16_port, 
      alu_out_s_15_port, alu_out_s_14_port, alu_out_s_13_port, 
      alu_out_s_12_port, alu_out_s_11_port, alu_out_s_10_port, alu_out_s_9_port
      , alu_out_s_8_port, alu_out_s_7_port, alu_out_s_6_port, alu_out_s_5_port,
      alu_out_s_4_port, alu_out_s_3_port, alu_out_s_2_port, alu_out_s_1_port, 
      alu_out_s_0_port, n17 : std_logic;

begin
   ZERO <= ZERO_port;
   
   MUXA : mux21_NBIT32_6 port map( A(31) => A_REG(31), A(30) => A_REG(30), 
                           A(29) => A_REG(29), A(28) => A_REG(28), A(27) => 
                           A_REG(27), A(26) => A_REG(26), A(25) => A_REG(25), 
                           A(24) => A_REG(24), A(23) => A_REG(23), A(22) => 
                           A_REG(22), A(21) => A_REG(21), A(20) => A_REG(20), 
                           A(19) => A_REG(19), A(18) => A_REG(18), A(17) => 
                           A_REG(17), A(16) => A_REG(16), A(15) => A_REG(15), 
                           A(14) => A_REG(14), A(13) => A_REG(13), A(12) => 
                           A_REG(12), A(11) => A_REG(11), A(10) => A_REG(10), 
                           A(9) => A_REG(9), A(8) => A_REG(8), A(7) => A_REG(7)
                           , A(6) => A_REG(6), A(5) => A_REG(5), A(4) => 
                           A_REG(4), A(3) => A_REG(3), A(2) => A_REG(2), A(1) 
                           => A_REG(1), A(0) => A_REG(0), B(31) => NPC_REG(31),
                           B(30) => NPC_REG(30), B(29) => NPC_REG(29), B(28) =>
                           NPC_REG(28), B(27) => NPC_REG(27), B(26) => 
                           NPC_REG(26), B(25) => NPC_REG(25), B(24) => 
                           NPC_REG(24), B(23) => NPC_REG(23), B(22) => 
                           NPC_REG(22), B(21) => NPC_REG(21), B(20) => 
                           NPC_REG(20), B(19) => NPC_REG(19), B(18) => 
                           NPC_REG(18), B(17) => NPC_REG(17), B(16) => 
                           NPC_REG(16), B(15) => NPC_REG(15), B(14) => 
                           NPC_REG(14), B(13) => NPC_REG(13), B(12) => 
                           NPC_REG(12), B(11) => NPC_REG(11), B(10) => 
                           NPC_REG(10), B(9) => NPC_REG(9), B(8) => NPC_REG(8),
                           B(7) => NPC_REG(7), B(6) => NPC_REG(6), B(5) => 
                           NPC_REG(5), B(4) => NPC_REG(4), B(3) => NPC_REG(3), 
                           B(2) => NPC_REG(2), B(1) => NPC_REG(1), B(0) => 
                           NPC_REG(0), sel => MUXA_SEL, muxout(31) => 
                           op_1_s_31_port, muxout(30) => op_1_s_30_port, 
                           muxout(29) => op_1_s_29_port, muxout(28) => 
                           op_1_s_28_port, muxout(27) => op_1_s_27_port, 
                           muxout(26) => op_1_s_26_port, muxout(25) => 
                           op_1_s_25_port, muxout(24) => op_1_s_24_port, 
                           muxout(23) => op_1_s_23_port, muxout(22) => 
                           op_1_s_22_port, muxout(21) => op_1_s_21_port, 
                           muxout(20) => op_1_s_20_port, muxout(19) => 
                           op_1_s_19_port, muxout(18) => op_1_s_18_port, 
                           muxout(17) => op_1_s_17_port, muxout(16) => 
                           op_1_s_16_port, muxout(15) => op_1_s_15_port, 
                           muxout(14) => op_1_s_14_port, muxout(13) => 
                           op_1_s_13_port, muxout(12) => op_1_s_12_port, 
                           muxout(11) => op_1_s_11_port, muxout(10) => 
                           op_1_s_10_port, muxout(9) => op_1_s_9_port, 
                           muxout(8) => op_1_s_8_port, muxout(7) => 
                           op_1_s_7_port, muxout(6) => op_1_s_6_port, muxout(5)
                           => op_1_s_5_port, muxout(4) => op_1_s_4_port, 
                           muxout(3) => op_1_s_3_port, muxout(2) => 
                           op_1_s_2_port, muxout(1) => op_1_s_1_port, muxout(0)
                           => op_1_s_0_port);
   MUXB : mux21_NBIT32_5 port map( A(31) => B_REG(31), A(30) => B_REG(30), 
                           A(29) => B_REG(29), A(28) => B_REG(28), A(27) => 
                           B_REG(27), A(26) => B_REG(26), A(25) => B_REG(25), 
                           A(24) => B_REG(24), A(23) => B_REG(23), A(22) => 
                           B_REG(22), A(21) => B_REG(21), A(20) => B_REG(20), 
                           A(19) => B_REG(19), A(18) => B_REG(18), A(17) => 
                           B_REG(17), A(16) => B_REG(16), A(15) => B_REG(15), 
                           A(14) => B_REG(14), A(13) => B_REG(13), A(12) => 
                           B_REG(12), A(11) => B_REG(11), A(10) => B_REG(10), 
                           A(9) => B_REG(9), A(8) => B_REG(8), A(7) => B_REG(7)
                           , A(6) => B_REG(6), A(5) => B_REG(5), A(4) => 
                           B_REG(4), A(3) => B_REG(3), A(2) => B_REG(2), A(1) 
                           => B_REG(1), A(0) => B_REG(0), B(31) => IMM_REG(31),
                           B(30) => IMM_REG(30), B(29) => IMM_REG(29), B(28) =>
                           IMM_REG(28), B(27) => IMM_REG(27), B(26) => 
                           IMM_REG(26), B(25) => IMM_REG(25), B(24) => 
                           IMM_REG(24), B(23) => IMM_REG(23), B(22) => 
                           IMM_REG(22), B(21) => IMM_REG(21), B(20) => 
                           IMM_REG(20), B(19) => IMM_REG(19), B(18) => 
                           IMM_REG(18), B(17) => IMM_REG(17), B(16) => 
                           IMM_REG(16), B(15) => IMM_REG(15), B(14) => 
                           IMM_REG(14), B(13) => IMM_REG(13), B(12) => 
                           IMM_REG(12), B(11) => IMM_REG(11), B(10) => 
                           IMM_REG(10), B(9) => IMM_REG(9), B(8) => IMM_REG(8),
                           B(7) => IMM_REG(7), B(6) => IMM_REG(6), B(5) => 
                           IMM_REG(5), B(4) => IMM_REG(4), B(3) => IMM_REG(3), 
                           B(2) => IMM_REG(2), B(1) => IMM_REG(1), B(0) => 
                           IMM_REG(0), sel => MUXB_SEL, muxout(31) => 
                           op_2_s_31_port, muxout(30) => op_2_s_30_port, 
                           muxout(29) => op_2_s_29_port, muxout(28) => 
                           op_2_s_28_port, muxout(27) => op_2_s_27_port, 
                           muxout(26) => op_2_s_26_port, muxout(25) => 
                           op_2_s_25_port, muxout(24) => op_2_s_24_port, 
                           muxout(23) => op_2_s_23_port, muxout(22) => 
                           op_2_s_22_port, muxout(21) => op_2_s_21_port, 
                           muxout(20) => op_2_s_20_port, muxout(19) => 
                           op_2_s_19_port, muxout(18) => op_2_s_18_port, 
                           muxout(17) => op_2_s_17_port, muxout(16) => 
                           op_2_s_16_port, muxout(15) => op_2_s_15_port, 
                           muxout(14) => op_2_s_14_port, muxout(13) => 
                           op_2_s_13_port, muxout(12) => op_2_s_12_port, 
                           muxout(11) => op_2_s_11_port, muxout(10) => 
                           op_2_s_10_port, muxout(9) => op_2_s_9_port, 
                           muxout(8) => op_2_s_8_port, muxout(7) => 
                           op_2_s_7_port, muxout(6) => op_2_s_6_port, muxout(5)
                           => op_2_s_5_port, muxout(4) => op_2_s_4_port, 
                           muxout(3) => op_2_s_3_port, muxout(2) => 
                           op_2_s_2_port, muxout(1) => op_2_s_1_port, muxout(0)
                           => op_2_s_0_port);
   MUX3 : mux21_NBIT32_4 port map( A(31) => alu_out_s_31_port, A(30) => 
                           alu_out_s_30_port, A(29) => alu_out_s_29_port, A(28)
                           => alu_out_s_28_port, A(27) => alu_out_s_27_port, 
                           A(26) => alu_out_s_26_port, A(25) => 
                           alu_out_s_25_port, A(24) => alu_out_s_24_port, A(23)
                           => alu_out_s_23_port, A(22) => alu_out_s_22_port, 
                           A(21) => alu_out_s_21_port, A(20) => 
                           alu_out_s_20_port, A(19) => alu_out_s_19_port, A(18)
                           => alu_out_s_18_port, A(17) => alu_out_s_17_port, 
                           A(16) => alu_out_s_16_port, A(15) => 
                           alu_out_s_15_port, A(14) => alu_out_s_14_port, A(13)
                           => alu_out_s_13_port, A(12) => alu_out_s_12_port, 
                           A(11) => alu_out_s_11_port, A(10) => 
                           alu_out_s_10_port, A(9) => alu_out_s_9_port, A(8) =>
                           alu_out_s_8_port, A(7) => alu_out_s_7_port, A(6) => 
                           alu_out_s_6_port, A(5) => alu_out_s_5_port, A(4) => 
                           alu_out_s_4_port, A(3) => alu_out_s_3_port, A(2) => 
                           alu_out_s_2_port, A(1) => alu_out_s_1_port, A(0) => 
                           alu_out_s_0_port, B(31) => PC_4(31), B(30) => 
                           PC_4(30), B(29) => PC_4(29), B(28) => PC_4(28), 
                           B(27) => PC_4(27), B(26) => PC_4(26), B(25) => 
                           PC_4(25), B(24) => PC_4(24), B(23) => PC_4(23), 
                           B(22) => PC_4(22), B(21) => PC_4(21), B(20) => 
                           PC_4(20), B(19) => PC_4(19), B(18) => PC_4(18), 
                           B(17) => PC_4(17), B(16) => PC_4(16), B(15) => 
                           PC_4(15), B(14) => PC_4(14), B(13) => PC_4(13), 
                           B(12) => PC_4(12), B(11) => PC_4(11), B(10) => 
                           PC_4(10), B(9) => PC_4(9), B(8) => PC_4(8), B(7) => 
                           PC_4(7), B(6) => PC_4(6), B(5) => PC_4(5), B(4) => 
                           PC_4(4), B(3) => PC_4(3), B(2) => PC_4(2), B(1) => 
                           PC_4(1), B(0) => PC_4(0), sel => ZERO_port, 
                           muxout(31) => BRANC_ADDR(31), muxout(30) => 
                           BRANC_ADDR(30), muxout(29) => BRANC_ADDR(29), 
                           muxout(28) => BRANC_ADDR(28), muxout(27) => 
                           BRANC_ADDR(27), muxout(26) => BRANC_ADDR(26), 
                           muxout(25) => BRANC_ADDR(25), muxout(24) => 
                           BRANC_ADDR(24), muxout(23) => BRANC_ADDR(23), 
                           muxout(22) => BRANC_ADDR(22), muxout(21) => 
                           BRANC_ADDR(21), muxout(20) => BRANC_ADDR(20), 
                           muxout(19) => BRANC_ADDR(19), muxout(18) => 
                           BRANC_ADDR(18), muxout(17) => BRANC_ADDR(17), 
                           muxout(16) => BRANC_ADDR(16), muxout(15) => 
                           BRANC_ADDR(15), muxout(14) => BRANC_ADDR(14), 
                           muxout(13) => BRANC_ADDR(13), muxout(12) => 
                           BRANC_ADDR(12), muxout(11) => BRANC_ADDR(11), 
                           muxout(10) => BRANC_ADDR(10), muxout(9) => 
                           BRANC_ADDR(9), muxout(8) => BRANC_ADDR(8), muxout(7)
                           => BRANC_ADDR(7), muxout(6) => BRANC_ADDR(6), 
                           muxout(5) => BRANC_ADDR(5), muxout(4) => 
                           BRANC_ADDR(4), muxout(3) => BRANC_ADDR(3), muxout(2)
                           => BRANC_ADDR(2), muxout(1) => BRANC_ADDR(1), 
                           muxout(0) => BRANC_ADDR(0));
   EXU_ALU : ALU_N32 port map( FUNC(0) => ALU_FUNC(0), FUNC(1) => ALU_FUNC(1), 
                           FUNC(2) => ALU_FUNC(2), FUNC(3) => ALU_FUNC(3), 
                           DATA1(31) => op_1_s_31_port, DATA1(30) => 
                           op_1_s_30_port, DATA1(29) => op_1_s_29_port, 
                           DATA1(28) => op_1_s_28_port, DATA1(27) => 
                           op_1_s_27_port, DATA1(26) => op_1_s_26_port, 
                           DATA1(25) => op_1_s_25_port, DATA1(24) => 
                           op_1_s_24_port, DATA1(23) => op_1_s_23_port, 
                           DATA1(22) => op_1_s_22_port, DATA1(21) => 
                           op_1_s_21_port, DATA1(20) => op_1_s_20_port, 
                           DATA1(19) => op_1_s_19_port, DATA1(18) => 
                           op_1_s_18_port, DATA1(17) => op_1_s_17_port, 
                           DATA1(16) => op_1_s_16_port, DATA1(15) => 
                           op_1_s_15_port, DATA1(14) => op_1_s_14_port, 
                           DATA1(13) => op_1_s_13_port, DATA1(12) => 
                           op_1_s_12_port, DATA1(11) => op_1_s_11_port, 
                           DATA1(10) => op_1_s_10_port, DATA1(9) => 
                           op_1_s_9_port, DATA1(8) => op_1_s_8_port, DATA1(7) 
                           => op_1_s_7_port, DATA1(6) => op_1_s_6_port, 
                           DATA1(5) => op_1_s_5_port, DATA1(4) => op_1_s_4_port
                           , DATA1(3) => op_1_s_3_port, DATA1(2) => 
                           op_1_s_2_port, DATA1(1) => op_1_s_1_port, DATA1(0) 
                           => op_1_s_0_port, DATA2(31) => op_2_s_31_port, 
                           DATA2(30) => op_2_s_30_port, DATA2(29) => 
                           op_2_s_29_port, DATA2(28) => op_2_s_28_port, 
                           DATA2(27) => op_2_s_27_port, DATA2(26) => 
                           op_2_s_26_port, DATA2(25) => op_2_s_25_port, 
                           DATA2(24) => op_2_s_24_port, DATA2(23) => 
                           op_2_s_23_port, DATA2(22) => op_2_s_22_port, 
                           DATA2(21) => op_2_s_21_port, DATA2(20) => 
                           op_2_s_20_port, DATA2(19) => op_2_s_19_port, 
                           DATA2(18) => op_2_s_18_port, DATA2(17) => 
                           op_2_s_17_port, DATA2(16) => op_2_s_16_port, 
                           DATA2(15) => op_2_s_15_port, DATA2(14) => 
                           op_2_s_14_port, DATA2(13) => op_2_s_13_port, 
                           DATA2(12) => op_2_s_12_port, DATA2(11) => 
                           op_2_s_11_port, DATA2(10) => op_2_s_10_port, 
                           DATA2(9) => op_2_s_9_port, DATA2(8) => op_2_s_8_port
                           , DATA2(7) => op_2_s_7_port, DATA2(6) => 
                           op_2_s_6_port, DATA2(5) => op_2_s_5_port, DATA2(4) 
                           => op_2_s_4_port, DATA2(3) => op_2_s_3_port, 
                           DATA2(2) => op_2_s_2_port, DATA2(1) => op_2_s_1_port
                           , DATA2(0) => op_2_s_0_port, OUTALU(31) => 
                           alu_out_s_31_port, OUTALU(30) => alu_out_s_30_port, 
                           OUTALU(29) => alu_out_s_29_port, OUTALU(28) => 
                           alu_out_s_28_port, OUTALU(27) => alu_out_s_27_port, 
                           OUTALU(26) => alu_out_s_26_port, OUTALU(25) => 
                           alu_out_s_25_port, OUTALU(24) => alu_out_s_24_port, 
                           OUTALU(23) => alu_out_s_23_port, OUTALU(22) => 
                           alu_out_s_22_port, OUTALU(21) => alu_out_s_21_port, 
                           OUTALU(20) => alu_out_s_20_port, OUTALU(19) => 
                           alu_out_s_19_port, OUTALU(18) => alu_out_s_18_port, 
                           OUTALU(17) => alu_out_s_17_port, OUTALU(16) => 
                           alu_out_s_16_port, OUTALU(15) => alu_out_s_15_port, 
                           OUTALU(14) => alu_out_s_14_port, OUTALU(13) => 
                           alu_out_s_13_port, OUTALU(12) => alu_out_s_12_port, 
                           OUTALU(11) => alu_out_s_11_port, OUTALU(10) => 
                           alu_out_s_10_port, OUTALU(9) => alu_out_s_9_port, 
                           OUTALU(8) => alu_out_s_8_port, OUTALU(7) => 
                           alu_out_s_7_port, OUTALU(6) => alu_out_s_6_port, 
                           OUTALU(5) => alu_out_s_5_port, OUTALU(4) => 
                           alu_out_s_4_port, OUTALU(3) => alu_out_s_3_port, 
                           OUTALU(2) => alu_out_s_2_port, OUTALU(1) => 
                           alu_out_s_1_port, OUTALU(0) => alu_out_s_0_port);
   EXU_CMPZ : is_zero_NBIT32 port map( A(31) => A_REG(31), A(30) => A_REG(30), 
                           A(29) => A_REG(29), A(28) => A_REG(28), A(27) => 
                           A_REG(27), A(26) => A_REG(26), A(25) => A_REG(25), 
                           A(24) => A_REG(24), A(23) => A_REG(23), A(22) => 
                           A_REG(22), A(21) => A_REG(21), A(20) => A_REG(20), 
                           A(19) => A_REG(19), A(18) => A_REG(18), A(17) => 
                           A_REG(17), A(16) => A_REG(16), A(15) => A_REG(15), 
                           A(14) => A_REG(14), A(13) => A_REG(13), A(12) => 
                           A_REG(12), A(11) => A_REG(11), A(10) => A_REG(10), 
                           A(9) => A_REG(9), A(8) => A_REG(8), A(7) => A_REG(7)
                           , A(6) => A_REG(6), A(5) => A_REG(5), A(4) => 
                           A_REG(4), A(3) => A_REG(3), A(2) => A_REG(2), A(1) 
                           => A_REG(1), A(0) => A_REG(0), BEQZ_OR_BNEZ => 
                           ZERO_SEL, EN => ZERO_EN, res => ZERO_port);
   NPC_REG_3 : reg_N32_7 port map( clk => CLK, rst => RST, en => n17, A(31) => 
                           NPC_REG(31), A(30) => NPC_REG(30), A(29) => 
                           NPC_REG(29), A(28) => NPC_REG(28), A(27) => 
                           NPC_REG(27), A(26) => NPC_REG(26), A(25) => 
                           NPC_REG(25), A(24) => NPC_REG(24), A(23) => 
                           NPC_REG(23), A(22) => NPC_REG(22), A(21) => 
                           NPC_REG(21), A(20) => NPC_REG(20), A(19) => 
                           NPC_REG(19), A(18) => NPC_REG(18), A(17) => 
                           NPC_REG(17), A(16) => NPC_REG(16), A(15) => 
                           NPC_REG(15), A(14) => NPC_REG(14), A(13) => 
                           NPC_REG(13), A(12) => NPC_REG(12), A(11) => 
                           NPC_REG(11), A(10) => NPC_REG(10), A(9) => 
                           NPC_REG(9), A(8) => NPC_REG(8), A(7) => NPC_REG(7), 
                           A(6) => NPC_REG(6), A(5) => NPC_REG(5), A(4) => 
                           NPC_REG(4), A(3) => NPC_REG(3), A(2) => NPC_REG(2), 
                           A(1) => NPC_REG(1), A(0) => NPC_REG(0), Y(31) => 
                           NPC_OUT(31), Y(30) => NPC_OUT(30), Y(29) => 
                           NPC_OUT(29), Y(28) => NPC_OUT(28), Y(27) => 
                           NPC_OUT(27), Y(26) => NPC_OUT(26), Y(25) => 
                           NPC_OUT(25), Y(24) => NPC_OUT(24), Y(23) => 
                           NPC_OUT(23), Y(22) => NPC_OUT(22), Y(21) => 
                           NPC_OUT(21), Y(20) => NPC_OUT(20), Y(19) => 
                           NPC_OUT(19), Y(18) => NPC_OUT(18), Y(17) => 
                           NPC_OUT(17), Y(16) => NPC_OUT(16), Y(15) => 
                           NPC_OUT(15), Y(14) => NPC_OUT(14), Y(13) => 
                           NPC_OUT(13), Y(12) => NPC_OUT(12), Y(11) => 
                           NPC_OUT(11), Y(10) => NPC_OUT(10), Y(9) => 
                           NPC_OUT(9), Y(8) => NPC_OUT(8), Y(7) => NPC_OUT(7), 
                           Y(6) => NPC_OUT(6), Y(5) => NPC_OUT(5), Y(4) => 
                           NPC_OUT(4), Y(3) => NPC_OUT(3), Y(2) => NPC_OUT(2), 
                           Y(1) => NPC_OUT(1), Y(0) => NPC_OUT(0));
   ALU_OUT_REG : reg_N32_6 port map( clk => CLK, rst => RST, en => ALUOUT_EN, 
                           A(31) => alu_out_s_31_port, A(30) => 
                           alu_out_s_30_port, A(29) => alu_out_s_29_port, A(28)
                           => alu_out_s_28_port, A(27) => alu_out_s_27_port, 
                           A(26) => alu_out_s_26_port, A(25) => 
                           alu_out_s_25_port, A(24) => alu_out_s_24_port, A(23)
                           => alu_out_s_23_port, A(22) => alu_out_s_22_port, 
                           A(21) => alu_out_s_21_port, A(20) => 
                           alu_out_s_20_port, A(19) => alu_out_s_19_port, A(18)
                           => alu_out_s_18_port, A(17) => alu_out_s_17_port, 
                           A(16) => alu_out_s_16_port, A(15) => 
                           alu_out_s_15_port, A(14) => alu_out_s_14_port, A(13)
                           => alu_out_s_13_port, A(12) => alu_out_s_12_port, 
                           A(11) => alu_out_s_11_port, A(10) => 
                           alu_out_s_10_port, A(9) => alu_out_s_9_port, A(8) =>
                           alu_out_s_8_port, A(7) => alu_out_s_7_port, A(6) => 
                           alu_out_s_6_port, A(5) => alu_out_s_5_port, A(4) => 
                           alu_out_s_4_port, A(3) => alu_out_s_3_port, A(2) => 
                           alu_out_s_2_port, A(1) => alu_out_s_1_port, A(0) => 
                           alu_out_s_0_port, Y(31) => ALU_OUT(31), Y(30) => 
                           ALU_OUT(30), Y(29) => ALU_OUT(29), Y(28) => 
                           ALU_OUT(28), Y(27) => ALU_OUT(27), Y(26) => 
                           ALU_OUT(26), Y(25) => ALU_OUT(25), Y(24) => 
                           ALU_OUT(24), Y(23) => ALU_OUT(23), Y(22) => 
                           ALU_OUT(22), Y(21) => ALU_OUT(21), Y(20) => 
                           ALU_OUT(20), Y(19) => ALU_OUT(19), Y(18) => 
                           ALU_OUT(18), Y(17) => ALU_OUT(17), Y(16) => 
                           ALU_OUT(16), Y(15) => ALU_OUT(15), Y(14) => 
                           ALU_OUT(14), Y(13) => ALU_OUT(13), Y(12) => 
                           ALU_OUT(12), Y(11) => ALU_OUT(11), Y(10) => 
                           ALU_OUT(10), Y(9) => ALU_OUT(9), Y(8) => ALU_OUT(8),
                           Y(7) => ALU_OUT(7), Y(6) => ALU_OUT(6), Y(5) => 
                           ALU_OUT(5), Y(4) => ALU_OUT(4), Y(3) => ALU_OUT(3), 
                           Y(2) => ALU_OUT(2), Y(1) => ALU_OUT(1), Y(0) => 
                           ALU_OUT(0));
   RT_REG_2 : reg_N32_5 port map( clk => CLK, rst => RST, en => n17, A(31) => 
                           RT_REG(31), A(30) => RT_REG(30), A(29) => RT_REG(29)
                           , A(28) => RT_REG(28), A(27) => RT_REG(27), A(26) =>
                           RT_REG(26), A(25) => RT_REG(25), A(24) => RT_REG(24)
                           , A(23) => RT_REG(23), A(22) => RT_REG(22), A(21) =>
                           RT_REG(21), A(20) => RT_REG(20), A(19) => RT_REG(19)
                           , A(18) => RT_REG(18), A(17) => RT_REG(17), A(16) =>
                           RT_REG(16), A(15) => RT_REG(15), A(14) => RT_REG(14)
                           , A(13) => RT_REG(13), A(12) => RT_REG(12), A(11) =>
                           RT_REG(11), A(10) => RT_REG(10), A(9) => RT_REG(9), 
                           A(8) => RT_REG(8), A(7) => RT_REG(7), A(6) => 
                           RT_REG(6), A(5) => RT_REG(5), A(4) => RT_REG(4), 
                           A(3) => RT_REG(3), A(2) => RT_REG(2), A(1) => 
                           RT_REG(1), A(0) => RT_REG(0), Y(31) => 
                           RT_REG_OUT(31), Y(30) => RT_REG_OUT(30), Y(29) => 
                           RT_REG_OUT(29), Y(28) => RT_REG_OUT(28), Y(27) => 
                           RT_REG_OUT(27), Y(26) => RT_REG_OUT(26), Y(25) => 
                           RT_REG_OUT(25), Y(24) => RT_REG_OUT(24), Y(23) => 
                           RT_REG_OUT(23), Y(22) => RT_REG_OUT(22), Y(21) => 
                           RT_REG_OUT(21), Y(20) => RT_REG_OUT(20), Y(19) => 
                           RT_REG_OUT(19), Y(18) => RT_REG_OUT(18), Y(17) => 
                           RT_REG_OUT(17), Y(16) => RT_REG_OUT(16), Y(15) => 
                           RT_REG_OUT(15), Y(14) => RT_REG_OUT(14), Y(13) => 
                           RT_REG_OUT(13), Y(12) => RT_REG_OUT(12), Y(11) => 
                           RT_REG_OUT(11), Y(10) => RT_REG_OUT(10), Y(9) => 
                           RT_REG_OUT(9), Y(8) => RT_REG_OUT(8), Y(7) => 
                           RT_REG_OUT(7), Y(6) => RT_REG_OUT(6), Y(5) => 
                           RT_REG_OUT(5), Y(4) => RT_REG_OUT(4), Y(3) => 
                           RT_REG_OUT(3), Y(2) => RT_REG_OUT(2), Y(1) => 
                           RT_REG_OUT(1), Y(0) => RT_REG_OUT(0));
   n17 <= '1';

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DU_N32 is

   port( J_EN, WR_EN, A_EN, B_EN, IMM_EN, RT_EN, is_R_type, BR_EN, clk, rst : 
         in std_logic;  NPC_IN, IR, DATAIN, ADDR_IN, BTA_OR_NPC : in 
         std_logic_vector (31 downto 0);  A, B, IMM, RT_OUT, NPC_OUT, PC_NXT : 
         out std_logic_vector (31 downto 0));

end DU_N32;

architecture SYN_struct of DU_N32 is

   component reg_N32_8
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   component adder_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  res : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component sign_extend_NBIT26_NBIT_F32
      port( A : in std_logic_vector (25 downto 0);  res : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component AND2
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component IV
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component reg_N32_9
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic;  
            muxout : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_10
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_extend_NBIT16_NBIT_F32
      port( A : in std_logic_vector (15 downto 0);  res : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component reg_N32_11
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_12
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_file_NBIT32_NREG32_NADDR5
      port( clk, rst, wr_en : in std_logic;  add_rd1, add_rd2 : in 
            std_logic_vector (4 downto 0);  add_wr, datain : in 
            std_logic_vector (31 downto 0);  out2, out1 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   signal B_nxt_31_port, B_nxt_30_port, B_nxt_29_port, B_nxt_28_port, 
      B_nxt_27_port, B_nxt_26_port, B_nxt_25_port, B_nxt_24_port, B_nxt_23_port
      , B_nxt_22_port, B_nxt_21_port, B_nxt_20_port, B_nxt_19_port, 
      B_nxt_18_port, B_nxt_17_port, B_nxt_16_port, B_nxt_15_port, B_nxt_14_port
      , B_nxt_13_port, B_nxt_12_port, B_nxt_11_port, B_nxt_10_port, 
      B_nxt_9_port, B_nxt_8_port, B_nxt_7_port, B_nxt_6_port, B_nxt_5_port, 
      B_nxt_4_port, B_nxt_3_port, B_nxt_2_port, B_nxt_1_port, B_nxt_0_port, 
      A_nxt_31_port, A_nxt_30_port, A_nxt_29_port, A_nxt_28_port, A_nxt_27_port
      , A_nxt_26_port, A_nxt_25_port, A_nxt_24_port, A_nxt_23_port, 
      A_nxt_22_port, A_nxt_21_port, A_nxt_20_port, A_nxt_19_port, A_nxt_18_port
      , A_nxt_17_port, A_nxt_16_port, A_nxt_15_port, A_nxt_14_port, 
      A_nxt_13_port, A_nxt_12_port, A_nxt_11_port, A_nxt_10_port, A_nxt_9_port,
      A_nxt_8_port, A_nxt_7_port, A_nxt_6_port, A_nxt_5_port, A_nxt_4_port, 
      A_nxt_3_port, A_nxt_2_port, A_nxt_1_port, A_nxt_0_port, IMM_nxt_31_port, 
      IMM_nxt_30_port, IMM_nxt_29_port, IMM_nxt_28_port, IMM_nxt_27_port, 
      IMM_nxt_26_port, IMM_nxt_25_port, IMM_nxt_24_port, IMM_nxt_23_port, 
      IMM_nxt_22_port, IMM_nxt_21_port, IMM_nxt_20_port, IMM_nxt_19_port, 
      IMM_nxt_18_port, IMM_nxt_17_port, IMM_nxt_16_port, IMM_nxt_15_port, 
      IMM_nxt_14_port, IMM_nxt_13_port, IMM_nxt_12_port, IMM_nxt_11_port, 
      IMM_nxt_10_port, IMM_nxt_9_port, IMM_nxt_8_port, IMM_nxt_7_port, 
      IMM_nxt_6_port, IMM_nxt_5_port, IMM_nxt_4_port, IMM_nxt_3_port, 
      IMM_nxt_2_port, IMM_nxt_1_port, IMM_nxt_0_port, BR_EN_NEG, J_SEL, 
      J_OFFSET_31_port, J_OFFSET_30_port, J_OFFSET_29_port, J_OFFSET_28_port, 
      J_OFFSET_27_port, J_OFFSET_26_port, J_OFFSET_25_port, J_OFFSET_24_port, 
      J_OFFSET_23_port, J_OFFSET_22_port, J_OFFSET_21_port, J_OFFSET_20_port, 
      J_OFFSET_19_port, J_OFFSET_18_port, J_OFFSET_17_port, J_OFFSET_16_port, 
      J_OFFSET_15_port, J_OFFSET_14_port, J_OFFSET_13_port, J_OFFSET_12_port, 
      J_OFFSET_11_port, J_OFFSET_10_port, J_OFFSET_9_port, J_OFFSET_8_port, 
      J_OFFSET_7_port, J_OFFSET_6_port, J_OFFSET_5_port, J_OFFSET_4_port, 
      J_OFFSET_3_port, J_OFFSET_2_port, J_OFFSET_1_port, J_OFFSET_0_port, 
      JTA_31_port, JTA_30_port, JTA_29_port, JTA_28_port, JTA_27_port, 
      JTA_26_port, JTA_25_port, JTA_24_port, JTA_23_port, JTA_22_port, 
      JTA_21_port, JTA_20_port, JTA_19_port, JTA_18_port, JTA_17_port, 
      JTA_16_port, JTA_15_port, JTA_14_port, JTA_13_port, JTA_12_port, 
      JTA_11_port, JTA_10_port, JTA_9_port, JTA_8_port, JTA_7_port, JTA_6_port,
      JTA_5_port, JTA_4_port, JTA_3_port, JTA_2_port, JTA_1_port, JTA_0_port, 
      RT_nxt_9_port, RT_nxt_8_port, RT_nxt_7_port, RT_nxt_6_port, RT_nxt_5_port
      , RT_nxt_4_port, RT_nxt_3_port, RT_nxt_31_port, RT_nxt_30_port, 
      RT_nxt_2_port, RT_nxt_29_port, RT_nxt_28_port, RT_nxt_27_port, 
      RT_nxt_26_port, RT_nxt_25_port, RT_nxt_24_port, RT_nxt_23_port, 
      RT_nxt_22_port, RT_nxt_21_port, RT_nxt_20_port, RT_nxt_1_port, 
      RT_nxt_19_port, RT_nxt_18_port, RT_nxt_17_port, RT_nxt_16_port, 
      RT_nxt_15_port, RT_nxt_14_port, RT_nxt_13_port, RT_nxt_12_port, 
      RT_nxt_11_port, RT_nxt_10_port, RT_nxt_0_port, n29, n30 : std_logic;

begin
   
   RF_instance : reg_file_NBIT32_NREG32_NADDR5 port map( clk => clk, rst => rst
                           , wr_en => WR_EN, add_rd1(4) => IR(25), add_rd1(3) 
                           => IR(24), add_rd1(2) => IR(23), add_rd1(1) => 
                           IR(22), add_rd1(0) => IR(21), add_rd2(4) => IR(20), 
                           add_rd2(3) => IR(19), add_rd2(2) => IR(18), 
                           add_rd2(1) => IR(17), add_rd2(0) => IR(16), 
                           add_wr(31) => ADDR_IN(31), add_wr(30) => ADDR_IN(30)
                           , add_wr(29) => ADDR_IN(29), add_wr(28) => 
                           ADDR_IN(28), add_wr(27) => ADDR_IN(27), add_wr(26) 
                           => ADDR_IN(26), add_wr(25) => ADDR_IN(25), 
                           add_wr(24) => ADDR_IN(24), add_wr(23) => ADDR_IN(23)
                           , add_wr(22) => ADDR_IN(22), add_wr(21) => 
                           ADDR_IN(21), add_wr(20) => ADDR_IN(20), add_wr(19) 
                           => ADDR_IN(19), add_wr(18) => ADDR_IN(18), 
                           add_wr(17) => ADDR_IN(17), add_wr(16) => ADDR_IN(16)
                           , add_wr(15) => ADDR_IN(15), add_wr(14) => 
                           ADDR_IN(14), add_wr(13) => ADDR_IN(13), add_wr(12) 
                           => ADDR_IN(12), add_wr(11) => ADDR_IN(11), 
                           add_wr(10) => ADDR_IN(10), add_wr(9) => ADDR_IN(9), 
                           add_wr(8) => ADDR_IN(8), add_wr(7) => ADDR_IN(7), 
                           add_wr(6) => ADDR_IN(6), add_wr(5) => ADDR_IN(5), 
                           add_wr(4) => ADDR_IN(4), add_wr(3) => ADDR_IN(3), 
                           add_wr(2) => ADDR_IN(2), add_wr(1) => ADDR_IN(1), 
                           add_wr(0) => ADDR_IN(0), datain(31) => DATAIN(31), 
                           datain(30) => DATAIN(30), datain(29) => DATAIN(29), 
                           datain(28) => DATAIN(28), datain(27) => DATAIN(27), 
                           datain(26) => DATAIN(26), datain(25) => DATAIN(25), 
                           datain(24) => DATAIN(24), datain(23) => DATAIN(23), 
                           datain(22) => DATAIN(22), datain(21) => DATAIN(21), 
                           datain(20) => DATAIN(20), datain(19) => DATAIN(19), 
                           datain(18) => DATAIN(18), datain(17) => DATAIN(17), 
                           datain(16) => DATAIN(16), datain(15) => DATAIN(15), 
                           datain(14) => DATAIN(14), datain(13) => DATAIN(13), 
                           datain(12) => DATAIN(12), datain(11) => DATAIN(11), 
                           datain(10) => DATAIN(10), datain(9) => DATAIN(9), 
                           datain(8) => DATAIN(8), datain(7) => DATAIN(7), 
                           datain(6) => DATAIN(6), datain(5) => DATAIN(5), 
                           datain(4) => DATAIN(4), datain(3) => DATAIN(3), 
                           datain(2) => DATAIN(2), datain(1) => DATAIN(1), 
                           datain(0) => DATAIN(0), out2(31) => B_nxt_31_port, 
                           out2(30) => B_nxt_30_port, out2(29) => B_nxt_29_port
                           , out2(28) => B_nxt_28_port, out2(27) => 
                           B_nxt_27_port, out2(26) => B_nxt_26_port, out2(25) 
                           => B_nxt_25_port, out2(24) => B_nxt_24_port, 
                           out2(23) => B_nxt_23_port, out2(22) => B_nxt_22_port
                           , out2(21) => B_nxt_21_port, out2(20) => 
                           B_nxt_20_port, out2(19) => B_nxt_19_port, out2(18) 
                           => B_nxt_18_port, out2(17) => B_nxt_17_port, 
                           out2(16) => B_nxt_16_port, out2(15) => B_nxt_15_port
                           , out2(14) => B_nxt_14_port, out2(13) => 
                           B_nxt_13_port, out2(12) => B_nxt_12_port, out2(11) 
                           => B_nxt_11_port, out2(10) => B_nxt_10_port, out2(9)
                           => B_nxt_9_port, out2(8) => B_nxt_8_port, out2(7) =>
                           B_nxt_7_port, out2(6) => B_nxt_6_port, out2(5) => 
                           B_nxt_5_port, out2(4) => B_nxt_4_port, out2(3) => 
                           B_nxt_3_port, out2(2) => B_nxt_2_port, out2(1) => 
                           B_nxt_1_port, out2(0) => B_nxt_0_port, out1(31) => 
                           A_nxt_31_port, out1(30) => A_nxt_30_port, out1(29) 
                           => A_nxt_29_port, out1(28) => A_nxt_28_port, 
                           out1(27) => A_nxt_27_port, out1(26) => A_nxt_26_port
                           , out1(25) => A_nxt_25_port, out1(24) => 
                           A_nxt_24_port, out1(23) => A_nxt_23_port, out1(22) 
                           => A_nxt_22_port, out1(21) => A_nxt_21_port, 
                           out1(20) => A_nxt_20_port, out1(19) => A_nxt_19_port
                           , out1(18) => A_nxt_18_port, out1(17) => 
                           A_nxt_17_port, out1(16) => A_nxt_16_port, out1(15) 
                           => A_nxt_15_port, out1(14) => A_nxt_14_port, 
                           out1(13) => A_nxt_13_port, out1(12) => A_nxt_12_port
                           , out1(11) => A_nxt_11_port, out1(10) => 
                           A_nxt_10_port, out1(9) => A_nxt_9_port, out1(8) => 
                           A_nxt_8_port, out1(7) => A_nxt_7_port, out1(6) => 
                           A_nxt_6_port, out1(5) => A_nxt_5_port, out1(4) => 
                           A_nxt_4_port, out1(3) => A_nxt_3_port, out1(2) => 
                           A_nxt_2_port, out1(1) => A_nxt_1_port, out1(0) => 
                           A_nxt_0_port);
   A_reg : reg_N32_12 port map( clk => clk, rst => rst, en => A_EN, A(31) => 
                           A_nxt_31_port, A(30) => A_nxt_30_port, A(29) => 
                           A_nxt_29_port, A(28) => A_nxt_28_port, A(27) => 
                           A_nxt_27_port, A(26) => A_nxt_26_port, A(25) => 
                           A_nxt_25_port, A(24) => A_nxt_24_port, A(23) => 
                           A_nxt_23_port, A(22) => A_nxt_22_port, A(21) => 
                           A_nxt_21_port, A(20) => A_nxt_20_port, A(19) => 
                           A_nxt_19_port, A(18) => A_nxt_18_port, A(17) => 
                           A_nxt_17_port, A(16) => A_nxt_16_port, A(15) => 
                           A_nxt_15_port, A(14) => A_nxt_14_port, A(13) => 
                           A_nxt_13_port, A(12) => A_nxt_12_port, A(11) => 
                           A_nxt_11_port, A(10) => A_nxt_10_port, A(9) => 
                           A_nxt_9_port, A(8) => A_nxt_8_port, A(7) => 
                           A_nxt_7_port, A(6) => A_nxt_6_port, A(5) => 
                           A_nxt_5_port, A(4) => A_nxt_4_port, A(3) => 
                           A_nxt_3_port, A(2) => A_nxt_2_port, A(1) => 
                           A_nxt_1_port, A(0) => A_nxt_0_port, Y(31) => A(31), 
                           Y(30) => A(30), Y(29) => A(29), Y(28) => A(28), 
                           Y(27) => A(27), Y(26) => A(26), Y(25) => A(25), 
                           Y(24) => A(24), Y(23) => A(23), Y(22) => A(22), 
                           Y(21) => A(21), Y(20) => A(20), Y(19) => A(19), 
                           Y(18) => A(18), Y(17) => A(17), Y(16) => A(16), 
                           Y(15) => A(15), Y(14) => A(14), Y(13) => A(13), 
                           Y(12) => A(12), Y(11) => A(11), Y(10) => A(10), Y(9)
                           => A(9), Y(8) => A(8), Y(7) => A(7), Y(6) => A(6), 
                           Y(5) => A(5), Y(4) => A(4), Y(3) => A(3), Y(2) => 
                           A(2), Y(1) => A(1), Y(0) => A(0));
   B_reg : reg_N32_11 port map( clk => clk, rst => rst, en => B_EN, A(31) => 
                           B_nxt_31_port, A(30) => B_nxt_30_port, A(29) => 
                           B_nxt_29_port, A(28) => B_nxt_28_port, A(27) => 
                           B_nxt_27_port, A(26) => B_nxt_26_port, A(25) => 
                           B_nxt_25_port, A(24) => B_nxt_24_port, A(23) => 
                           B_nxt_23_port, A(22) => B_nxt_22_port, A(21) => 
                           B_nxt_21_port, A(20) => B_nxt_20_port, A(19) => 
                           B_nxt_19_port, A(18) => B_nxt_18_port, A(17) => 
                           B_nxt_17_port, A(16) => B_nxt_16_port, A(15) => 
                           B_nxt_15_port, A(14) => B_nxt_14_port, A(13) => 
                           B_nxt_13_port, A(12) => B_nxt_12_port, A(11) => 
                           B_nxt_11_port, A(10) => B_nxt_10_port, A(9) => 
                           B_nxt_9_port, A(8) => B_nxt_8_port, A(7) => 
                           B_nxt_7_port, A(6) => B_nxt_6_port, A(5) => 
                           B_nxt_5_port, A(4) => B_nxt_4_port, A(3) => 
                           B_nxt_3_port, A(2) => B_nxt_2_port, A(1) => 
                           B_nxt_1_port, A(0) => B_nxt_0_port, Y(31) => B(31), 
                           Y(30) => B(30), Y(29) => B(29), Y(28) => B(28), 
                           Y(27) => B(27), Y(26) => B(26), Y(25) => B(25), 
                           Y(24) => B(24), Y(23) => B(23), Y(22) => B(22), 
                           Y(21) => B(21), Y(20) => B(20), Y(19) => B(19), 
                           Y(18) => B(18), Y(17) => B(17), Y(16) => B(16), 
                           Y(15) => B(15), Y(14) => B(14), Y(13) => B(13), 
                           Y(12) => B(12), Y(11) => B(11), Y(10) => B(10), Y(9)
                           => B(9), Y(8) => B(8), Y(7) => B(7), Y(6) => B(6), 
                           Y(5) => B(5), Y(4) => B(4), Y(3) => B(3), Y(2) => 
                           B(2), Y(1) => B(1), Y(0) => B(0));
   Sign_extend_block : sign_extend_NBIT16_NBIT_F32 port map( A(15) => IR(15), 
                           A(14) => IR(14), A(13) => IR(13), A(12) => IR(12), 
                           A(11) => IR(11), A(10) => IR(10), A(9) => IR(9), 
                           A(8) => IR(8), A(7) => IR(7), A(6) => IR(6), A(5) =>
                           IR(5), A(4) => IR(4), A(3) => IR(3), A(2) => IR(2), 
                           A(1) => IR(1), A(0) => IR(0), res(31) => 
                           IMM_nxt_31_port, res(30) => IMM_nxt_30_port, res(29)
                           => IMM_nxt_29_port, res(28) => IMM_nxt_28_port, 
                           res(27) => IMM_nxt_27_port, res(26) => 
                           IMM_nxt_26_port, res(25) => IMM_nxt_25_port, res(24)
                           => IMM_nxt_24_port, res(23) => IMM_nxt_23_port, 
                           res(22) => IMM_nxt_22_port, res(21) => 
                           IMM_nxt_21_port, res(20) => IMM_nxt_20_port, res(19)
                           => IMM_nxt_19_port, res(18) => IMM_nxt_18_port, 
                           res(17) => IMM_nxt_17_port, res(16) => 
                           IMM_nxt_16_port, res(15) => IMM_nxt_15_port, res(14)
                           => IMM_nxt_14_port, res(13) => IMM_nxt_13_port, 
                           res(12) => IMM_nxt_12_port, res(11) => 
                           IMM_nxt_11_port, res(10) => IMM_nxt_10_port, res(9) 
                           => IMM_nxt_9_port, res(8) => IMM_nxt_8_port, res(7) 
                           => IMM_nxt_7_port, res(6) => IMM_nxt_6_port, res(5) 
                           => IMM_nxt_5_port, res(4) => IMM_nxt_4_port, res(3) 
                           => IMM_nxt_3_port, res(2) => IMM_nxt_2_port, res(1) 
                           => IMM_nxt_1_port, res(0) => IMM_nxt_0_port);
   IMM_reg : reg_N32_10 port map( clk => clk, rst => rst, en => IMM_EN, A(31) 
                           => IMM_nxt_31_port, A(30) => IMM_nxt_30_port, A(29) 
                           => IMM_nxt_29_port, A(28) => IMM_nxt_28_port, A(27) 
                           => IMM_nxt_27_port, A(26) => IMM_nxt_26_port, A(25) 
                           => IMM_nxt_25_port, A(24) => IMM_nxt_24_port, A(23) 
                           => IMM_nxt_23_port, A(22) => IMM_nxt_22_port, A(21) 
                           => IMM_nxt_21_port, A(20) => IMM_nxt_20_port, A(19) 
                           => IMM_nxt_19_port, A(18) => IMM_nxt_18_port, A(17) 
                           => IMM_nxt_17_port, A(16) => IMM_nxt_16_port, A(15) 
                           => IMM_nxt_15_port, A(14) => IMM_nxt_14_port, A(13) 
                           => IMM_nxt_13_port, A(12) => IMM_nxt_12_port, A(11) 
                           => IMM_nxt_11_port, A(10) => IMM_nxt_10_port, A(9) 
                           => IMM_nxt_9_port, A(8) => IMM_nxt_8_port, A(7) => 
                           IMM_nxt_7_port, A(6) => IMM_nxt_6_port, A(5) => 
                           IMM_nxt_5_port, A(4) => IMM_nxt_4_port, A(3) => 
                           IMM_nxt_3_port, A(2) => IMM_nxt_2_port, A(1) => 
                           IMM_nxt_1_port, A(0) => IMM_nxt_0_port, Y(31) => 
                           IMM(31), Y(30) => IMM(30), Y(29) => IMM(29), Y(28) 
                           => IMM(28), Y(27) => IMM(27), Y(26) => IMM(26), 
                           Y(25) => IMM(25), Y(24) => IMM(24), Y(23) => IMM(23)
                           , Y(22) => IMM(22), Y(21) => IMM(21), Y(20) => 
                           IMM(20), Y(19) => IMM(19), Y(18) => IMM(18), Y(17) 
                           => IMM(17), Y(16) => IMM(16), Y(15) => IMM(15), 
                           Y(14) => IMM(14), Y(13) => IMM(13), Y(12) => IMM(12)
                           , Y(11) => IMM(11), Y(10) => IMM(10), Y(9) => IMM(9)
                           , Y(8) => IMM(8), Y(7) => IMM(7), Y(6) => IMM(6), 
                           Y(5) => IMM(5), Y(4) => IMM(4), Y(3) => IMM(3), Y(2)
                           => IMM(2), Y(1) => IMM(1), Y(0) => IMM(0));
   RT_source_mux : mux21_NBIT32_0 port map( A(31) => n30, A(30) => n30, A(29) 
                           => n30, A(28) => n30, A(27) => n30, A(26) => n30, 
                           A(25) => n30, A(24) => n30, A(23) => n30, A(22) => 
                           n30, A(21) => n30, A(20) => n30, A(19) => n30, A(18)
                           => n30, A(17) => n30, A(16) => n30, A(15) => n30, 
                           A(14) => n30, A(13) => n30, A(12) => n30, A(11) => 
                           n30, A(10) => n30, A(9) => n30, A(8) => n30, A(7) =>
                           n30, A(6) => n30, A(5) => n30, A(4) => IR(15), A(3) 
                           => IR(14), A(2) => IR(13), A(1) => IR(12), A(0) => 
                           IR(11), B(31) => n30, B(30) => n30, B(29) => n30, 
                           B(28) => n30, B(27) => n30, B(26) => n30, B(25) => 
                           n30, B(24) => n30, B(23) => n30, B(22) => n30, B(21)
                           => n30, B(20) => n30, B(19) => n30, B(18) => n30, 
                           B(17) => n30, B(16) => n30, B(15) => n30, B(14) => 
                           n30, B(13) => n30, B(12) => n30, B(11) => n30, B(10)
                           => n30, B(9) => n30, B(8) => n30, B(7) => n30, B(6) 
                           => n30, B(5) => n30, B(4) => IR(20), B(3) => IR(19),
                           B(2) => IR(18), B(1) => IR(17), B(0) => IR(16), sel 
                           => is_R_type, muxout(31) => RT_nxt_31_port, 
                           muxout(30) => RT_nxt_30_port, muxout(29) => 
                           RT_nxt_29_port, muxout(28) => RT_nxt_28_port, 
                           muxout(27) => RT_nxt_27_port, muxout(26) => 
                           RT_nxt_26_port, muxout(25) => RT_nxt_25_port, 
                           muxout(24) => RT_nxt_24_port, muxout(23) => 
                           RT_nxt_23_port, muxout(22) => RT_nxt_22_port, 
                           muxout(21) => RT_nxt_21_port, muxout(20) => 
                           RT_nxt_20_port, muxout(19) => RT_nxt_19_port, 
                           muxout(18) => RT_nxt_18_port, muxout(17) => 
                           RT_nxt_17_port, muxout(16) => RT_nxt_16_port, 
                           muxout(15) => RT_nxt_15_port, muxout(14) => 
                           RT_nxt_14_port, muxout(13) => RT_nxt_13_port, 
                           muxout(12) => RT_nxt_12_port, muxout(11) => 
                           RT_nxt_11_port, muxout(10) => RT_nxt_10_port, 
                           muxout(9) => RT_nxt_9_port, muxout(8) => 
                           RT_nxt_8_port, muxout(7) => RT_nxt_7_port, muxout(6)
                           => RT_nxt_6_port, muxout(5) => RT_nxt_5_port, 
                           muxout(4) => RT_nxt_4_port, muxout(3) => 
                           RT_nxt_3_port, muxout(2) => RT_nxt_2_port, muxout(1)
                           => RT_nxt_1_port, muxout(0) => RT_nxt_0_port);
   RT_reg_inst : reg_N32_9 port map( clk => clk, rst => rst, en => RT_EN, A(31)
                           => RT_nxt_31_port, A(30) => RT_nxt_30_port, A(29) =>
                           RT_nxt_29_port, A(28) => RT_nxt_28_port, A(27) => 
                           RT_nxt_27_port, A(26) => RT_nxt_26_port, A(25) => 
                           RT_nxt_25_port, A(24) => RT_nxt_24_port, A(23) => 
                           RT_nxt_23_port, A(22) => RT_nxt_22_port, A(21) => 
                           RT_nxt_21_port, A(20) => RT_nxt_20_port, A(19) => 
                           RT_nxt_19_port, A(18) => RT_nxt_18_port, A(17) => 
                           RT_nxt_17_port, A(16) => RT_nxt_16_port, A(15) => 
                           RT_nxt_15_port, A(14) => RT_nxt_14_port, A(13) => 
                           RT_nxt_13_port, A(12) => RT_nxt_12_port, A(11) => 
                           RT_nxt_11_port, A(10) => RT_nxt_10_port, A(9) => 
                           RT_nxt_9_port, A(8) => RT_nxt_8_port, A(7) => 
                           RT_nxt_7_port, A(6) => RT_nxt_6_port, A(5) => 
                           RT_nxt_5_port, A(4) => RT_nxt_4_port, A(3) => 
                           RT_nxt_3_port, A(2) => RT_nxt_2_port, A(1) => 
                           RT_nxt_1_port, A(0) => RT_nxt_0_port, Y(31) => 
                           RT_OUT(31), Y(30) => RT_OUT(30), Y(29) => RT_OUT(29)
                           , Y(28) => RT_OUT(28), Y(27) => RT_OUT(27), Y(26) =>
                           RT_OUT(26), Y(25) => RT_OUT(25), Y(24) => RT_OUT(24)
                           , Y(23) => RT_OUT(23), Y(22) => RT_OUT(22), Y(21) =>
                           RT_OUT(21), Y(20) => RT_OUT(20), Y(19) => RT_OUT(19)
                           , Y(18) => RT_OUT(18), Y(17) => RT_OUT(17), Y(16) =>
                           RT_OUT(16), Y(15) => RT_OUT(15), Y(14) => RT_OUT(14)
                           , Y(13) => RT_OUT(13), Y(12) => RT_OUT(12), Y(11) =>
                           RT_OUT(11), Y(10) => RT_OUT(10), Y(9) => RT_OUT(9), 
                           Y(8) => RT_OUT(8), Y(7) => RT_OUT(7), Y(6) => 
                           RT_OUT(6), Y(5) => RT_OUT(5), Y(4) => RT_OUT(4), 
                           Y(3) => RT_OUT(3), Y(2) => RT_OUT(2), Y(1) => 
                           RT_OUT(1), Y(0) => RT_OUT(0));
   IV_instance : IV port map( A => BR_EN, Y => BR_EN_NEG);
   AND2_instance : AND2 port map( a => BR_EN_NEG, b => J_EN, y => J_SEL);
   addr_sign_extend : sign_extend_NBIT26_NBIT_F32 port map( A(25) => IR(25), 
                           A(24) => IR(24), A(23) => IR(23), A(22) => IR(22), 
                           A(21) => IR(21), A(20) => IR(20), A(19) => IR(19), 
                           A(18) => IR(18), A(17) => IR(17), A(16) => IR(16), 
                           A(15) => IR(15), A(14) => IR(14), A(13) => IR(13), 
                           A(12) => IR(12), A(11) => IR(11), A(10) => IR(10), 
                           A(9) => IR(9), A(8) => IR(8), A(7) => IR(7), A(6) =>
                           IR(6), A(5) => IR(5), A(4) => IR(4), A(3) => IR(3), 
                           A(2) => IR(2), A(1) => IR(1), A(0) => IR(0), res(31)
                           => J_OFFSET_31_port, res(30) => J_OFFSET_30_port, 
                           res(29) => J_OFFSET_29_port, res(28) => 
                           J_OFFSET_28_port, res(27) => J_OFFSET_27_port, 
                           res(26) => J_OFFSET_26_port, res(25) => 
                           J_OFFSET_25_port, res(24) => J_OFFSET_24_port, 
                           res(23) => J_OFFSET_23_port, res(22) => 
                           J_OFFSET_22_port, res(21) => J_OFFSET_21_port, 
                           res(20) => J_OFFSET_20_port, res(19) => 
                           J_OFFSET_19_port, res(18) => J_OFFSET_18_port, 
                           res(17) => J_OFFSET_17_port, res(16) => 
                           J_OFFSET_16_port, res(15) => J_OFFSET_15_port, 
                           res(14) => J_OFFSET_14_port, res(13) => 
                           J_OFFSET_13_port, res(12) => J_OFFSET_12_port, 
                           res(11) => J_OFFSET_11_port, res(10) => 
                           J_OFFSET_10_port, res(9) => J_OFFSET_9_port, res(8) 
                           => J_OFFSET_8_port, res(7) => J_OFFSET_7_port, 
                           res(6) => J_OFFSET_6_port, res(5) => J_OFFSET_5_port
                           , res(4) => J_OFFSET_4_port, res(3) => 
                           J_OFFSET_3_port, res(2) => J_OFFSET_2_port, res(1) 
                           => J_OFFSET_1_port, res(0) => J_OFFSET_0_port);
   ADD_instance : adder_NBIT32 port map( A(31) => NPC_IN(31), A(30) => 
                           NPC_IN(30), A(29) => NPC_IN(29), A(28) => NPC_IN(28)
                           , A(27) => NPC_IN(27), A(26) => NPC_IN(26), A(25) =>
                           NPC_IN(25), A(24) => NPC_IN(24), A(23) => NPC_IN(23)
                           , A(22) => NPC_IN(22), A(21) => NPC_IN(21), A(20) =>
                           NPC_IN(20), A(19) => NPC_IN(19), A(18) => NPC_IN(18)
                           , A(17) => NPC_IN(17), A(16) => NPC_IN(16), A(15) =>
                           NPC_IN(15), A(14) => NPC_IN(14), A(13) => NPC_IN(13)
                           , A(12) => NPC_IN(12), A(11) => NPC_IN(11), A(10) =>
                           NPC_IN(10), A(9) => NPC_IN(9), A(8) => NPC_IN(8), 
                           A(7) => NPC_IN(7), A(6) => NPC_IN(6), A(5) => 
                           NPC_IN(5), A(4) => NPC_IN(4), A(3) => NPC_IN(3), 
                           A(2) => NPC_IN(2), A(1) => NPC_IN(1), A(0) => 
                           NPC_IN(0), B(31) => J_OFFSET_31_port, B(30) => 
                           J_OFFSET_30_port, B(29) => J_OFFSET_29_port, B(28) 
                           => J_OFFSET_28_port, B(27) => J_OFFSET_27_port, 
                           B(26) => J_OFFSET_26_port, B(25) => J_OFFSET_25_port
                           , B(24) => J_OFFSET_24_port, B(23) => 
                           J_OFFSET_23_port, B(22) => J_OFFSET_22_port, B(21) 
                           => J_OFFSET_21_port, B(20) => J_OFFSET_20_port, 
                           B(19) => J_OFFSET_19_port, B(18) => J_OFFSET_18_port
                           , B(17) => J_OFFSET_17_port, B(16) => 
                           J_OFFSET_16_port, B(15) => J_OFFSET_15_port, B(14) 
                           => J_OFFSET_14_port, B(13) => J_OFFSET_13_port, 
                           B(12) => J_OFFSET_12_port, B(11) => J_OFFSET_11_port
                           , B(10) => J_OFFSET_10_port, B(9) => J_OFFSET_9_port
                           , B(8) => J_OFFSET_8_port, B(7) => J_OFFSET_7_port, 
                           B(6) => J_OFFSET_6_port, B(5) => J_OFFSET_5_port, 
                           B(4) => J_OFFSET_4_port, B(3) => J_OFFSET_3_port, 
                           B(2) => J_OFFSET_2_port, B(1) => J_OFFSET_1_port, 
                           B(0) => J_OFFSET_0_port, res(31) => JTA_31_port, 
                           res(30) => JTA_30_port, res(29) => JTA_29_port, 
                           res(28) => JTA_28_port, res(27) => JTA_27_port, 
                           res(26) => JTA_26_port, res(25) => JTA_25_port, 
                           res(24) => JTA_24_port, res(23) => JTA_23_port, 
                           res(22) => JTA_22_port, res(21) => JTA_21_port, 
                           res(20) => JTA_20_port, res(19) => JTA_19_port, 
                           res(18) => JTA_18_port, res(17) => JTA_17_port, 
                           res(16) => JTA_16_port, res(15) => JTA_15_port, 
                           res(14) => JTA_14_port, res(13) => JTA_13_port, 
                           res(12) => JTA_12_port, res(11) => JTA_11_port, 
                           res(10) => JTA_10_port, res(9) => JTA_9_port, res(8)
                           => JTA_8_port, res(7) => JTA_7_port, res(6) => 
                           JTA_6_port, res(5) => JTA_5_port, res(4) => 
                           JTA_4_port, res(3) => JTA_3_port, res(2) => 
                           JTA_2_port, res(1) => JTA_1_port, res(0) => 
                           JTA_0_port);
   PC_source_MUX : mux21_NBIT32_7 port map( A(31) => JTA_31_port, A(30) => 
                           JTA_30_port, A(29) => JTA_29_port, A(28) => 
                           JTA_28_port, A(27) => JTA_27_port, A(26) => 
                           JTA_26_port, A(25) => JTA_25_port, A(24) => 
                           JTA_24_port, A(23) => JTA_23_port, A(22) => 
                           JTA_22_port, A(21) => JTA_21_port, A(20) => 
                           JTA_20_port, A(19) => JTA_19_port, A(18) => 
                           JTA_18_port, A(17) => JTA_17_port, A(16) => 
                           JTA_16_port, A(15) => JTA_15_port, A(14) => 
                           JTA_14_port, A(13) => JTA_13_port, A(12) => 
                           JTA_12_port, A(11) => JTA_11_port, A(10) => 
                           JTA_10_port, A(9) => JTA_9_port, A(8) => JTA_8_port,
                           A(7) => JTA_7_port, A(6) => JTA_6_port, A(5) => 
                           JTA_5_port, A(4) => JTA_4_port, A(3) => JTA_3_port, 
                           A(2) => JTA_2_port, A(1) => JTA_1_port, A(0) => 
                           JTA_0_port, B(31) => BTA_OR_NPC(31), B(30) => 
                           BTA_OR_NPC(30), B(29) => BTA_OR_NPC(29), B(28) => 
                           BTA_OR_NPC(28), B(27) => BTA_OR_NPC(27), B(26) => 
                           BTA_OR_NPC(26), B(25) => BTA_OR_NPC(25), B(24) => 
                           BTA_OR_NPC(24), B(23) => BTA_OR_NPC(23), B(22) => 
                           BTA_OR_NPC(22), B(21) => BTA_OR_NPC(21), B(20) => 
                           BTA_OR_NPC(20), B(19) => BTA_OR_NPC(19), B(18) => 
                           BTA_OR_NPC(18), B(17) => BTA_OR_NPC(17), B(16) => 
                           BTA_OR_NPC(16), B(15) => BTA_OR_NPC(15), B(14) => 
                           BTA_OR_NPC(14), B(13) => BTA_OR_NPC(13), B(12) => 
                           BTA_OR_NPC(12), B(11) => BTA_OR_NPC(11), B(10) => 
                           BTA_OR_NPC(10), B(9) => BTA_OR_NPC(9), B(8) => 
                           BTA_OR_NPC(8), B(7) => BTA_OR_NPC(7), B(6) => 
                           BTA_OR_NPC(6), B(5) => BTA_OR_NPC(5), B(4) => 
                           BTA_OR_NPC(4), B(3) => BTA_OR_NPC(3), B(2) => 
                           BTA_OR_NPC(2), B(1) => BTA_OR_NPC(1), B(0) => 
                           BTA_OR_NPC(0), sel => J_SEL, muxout(31) => 
                           PC_NXT(31), muxout(30) => PC_NXT(30), muxout(29) => 
                           PC_NXT(29), muxout(28) => PC_NXT(28), muxout(27) => 
                           PC_NXT(27), muxout(26) => PC_NXT(26), muxout(25) => 
                           PC_NXT(25), muxout(24) => PC_NXT(24), muxout(23) => 
                           PC_NXT(23), muxout(22) => PC_NXT(22), muxout(21) => 
                           PC_NXT(21), muxout(20) => PC_NXT(20), muxout(19) => 
                           PC_NXT(19), muxout(18) => PC_NXT(18), muxout(17) => 
                           PC_NXT(17), muxout(16) => PC_NXT(16), muxout(15) => 
                           PC_NXT(15), muxout(14) => PC_NXT(14), muxout(13) => 
                           PC_NXT(13), muxout(12) => PC_NXT(12), muxout(11) => 
                           PC_NXT(11), muxout(10) => PC_NXT(10), muxout(9) => 
                           PC_NXT(9), muxout(8) => PC_NXT(8), muxout(7) => 
                           PC_NXT(7), muxout(6) => PC_NXT(6), muxout(5) => 
                           PC_NXT(5), muxout(4) => PC_NXT(4), muxout(3) => 
                           PC_NXT(3), muxout(2) => PC_NXT(2), muxout(1) => 
                           PC_NXT(1), muxout(0) => PC_NXT(0));
   NPC_reg_inst : reg_N32_8 port map( clk => clk, rst => rst, en => n29, A(31) 
                           => NPC_IN(31), A(30) => NPC_IN(30), A(29) => 
                           NPC_IN(29), A(28) => NPC_IN(28), A(27) => NPC_IN(27)
                           , A(26) => NPC_IN(26), A(25) => NPC_IN(25), A(24) =>
                           NPC_IN(24), A(23) => NPC_IN(23), A(22) => NPC_IN(22)
                           , A(21) => NPC_IN(21), A(20) => NPC_IN(20), A(19) =>
                           NPC_IN(19), A(18) => NPC_IN(18), A(17) => NPC_IN(17)
                           , A(16) => NPC_IN(16), A(15) => NPC_IN(15), A(14) =>
                           NPC_IN(14), A(13) => NPC_IN(13), A(12) => NPC_IN(12)
                           , A(11) => NPC_IN(11), A(10) => NPC_IN(10), A(9) => 
                           NPC_IN(9), A(8) => NPC_IN(8), A(7) => NPC_IN(7), 
                           A(6) => NPC_IN(6), A(5) => NPC_IN(5), A(4) => 
                           NPC_IN(4), A(3) => NPC_IN(3), A(2) => NPC_IN(2), 
                           A(1) => NPC_IN(1), A(0) => NPC_IN(0), Y(31) => 
                           NPC_OUT(31), Y(30) => NPC_OUT(30), Y(29) => 
                           NPC_OUT(29), Y(28) => NPC_OUT(28), Y(27) => 
                           NPC_OUT(27), Y(26) => NPC_OUT(26), Y(25) => 
                           NPC_OUT(25), Y(24) => NPC_OUT(24), Y(23) => 
                           NPC_OUT(23), Y(22) => NPC_OUT(22), Y(21) => 
                           NPC_OUT(21), Y(20) => NPC_OUT(20), Y(19) => 
                           NPC_OUT(19), Y(18) => NPC_OUT(18), Y(17) => 
                           NPC_OUT(17), Y(16) => NPC_OUT(16), Y(15) => 
                           NPC_OUT(15), Y(14) => NPC_OUT(14), Y(13) => 
                           NPC_OUT(13), Y(12) => NPC_OUT(12), Y(11) => 
                           NPC_OUT(11), Y(10) => NPC_OUT(10), Y(9) => 
                           NPC_OUT(9), Y(8) => NPC_OUT(8), Y(7) => NPC_OUT(7), 
                           Y(6) => NPC_OUT(6), Y(5) => NPC_OUT(5), Y(4) => 
                           NPC_OUT(4), Y(3) => NPC_OUT(3), Y(2) => NPC_OUT(2), 
                           Y(1) => NPC_OUT(1), Y(0) => NPC_OUT(0));
   n29 <= '1';
   n30 <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FU_N32 is

   port( CLK, RST, PC_EN, NPC_EN, IR_EN : in std_logic;  IN_ID, from_IRAM : in 
         std_logic_vector (31 downto 0);  to_IRAM, IREG_out, NPC_out, PC_4out :
         out std_logic_vector (31 downto 0));

end FU_N32;

architecture SYN_structural of FU_N32 is

   component reg_N32_13
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_N32_14
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component add4_NBIT32
      port( A : in std_logic_vector (31 downto 0);  res : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component reg_N32_0
      port( clk, rst, en : in std_logic;  A : in std_logic_vector (31 downto 0)
            ;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   signal to_IRAM_31_port, to_IRAM_30_port, to_IRAM_29_port, to_IRAM_28_port, 
      to_IRAM_27_port, to_IRAM_26_port, to_IRAM_25_port, to_IRAM_24_port, 
      to_IRAM_23_port, to_IRAM_22_port, to_IRAM_21_port, to_IRAM_20_port, 
      to_IRAM_19_port, to_IRAM_18_port, to_IRAM_17_port, to_IRAM_16_port, 
      to_IRAM_15_port, to_IRAM_14_port, to_IRAM_13_port, to_IRAM_12_port, 
      to_IRAM_11_port, to_IRAM_10_port, to_IRAM_9_port, to_IRAM_8_port, 
      to_IRAM_7_port, to_IRAM_6_port, to_IRAM_5_port, to_IRAM_4_port, 
      to_IRAM_3_port, to_IRAM_2_port, to_IRAM_1_port, to_IRAM_0_port, 
      PC_4out_31_port, PC_4out_30_port, PC_4out_29_port, PC_4out_28_port, 
      PC_4out_27_port, PC_4out_26_port, PC_4out_25_port, PC_4out_24_port, 
      PC_4out_23_port, PC_4out_22_port, PC_4out_21_port, PC_4out_20_port, 
      PC_4out_19_port, PC_4out_18_port, PC_4out_17_port, PC_4out_16_port, 
      PC_4out_15_port, PC_4out_14_port, PC_4out_13_port, PC_4out_12_port, 
      PC_4out_11_port, PC_4out_10_port, PC_4out_9_port, PC_4out_8_port, 
      PC_4out_7_port, PC_4out_6_port, PC_4out_5_port, PC_4out_4_port, 
      PC_4out_3_port, PC_4out_2_port, PC_4out_1_port, PC_4out_0_port : 
      std_logic;

begin
   to_IRAM <= ( to_IRAM_31_port, to_IRAM_30_port, to_IRAM_29_port, 
      to_IRAM_28_port, to_IRAM_27_port, to_IRAM_26_port, to_IRAM_25_port, 
      to_IRAM_24_port, to_IRAM_23_port, to_IRAM_22_port, to_IRAM_21_port, 
      to_IRAM_20_port, to_IRAM_19_port, to_IRAM_18_port, to_IRAM_17_port, 
      to_IRAM_16_port, to_IRAM_15_port, to_IRAM_14_port, to_IRAM_13_port, 
      to_IRAM_12_port, to_IRAM_11_port, to_IRAM_10_port, to_IRAM_9_port, 
      to_IRAM_8_port, to_IRAM_7_port, to_IRAM_6_port, to_IRAM_5_port, 
      to_IRAM_4_port, to_IRAM_3_port, to_IRAM_2_port, to_IRAM_1_port, 
      to_IRAM_0_port );
   PC_4out <= ( PC_4out_31_port, PC_4out_30_port, PC_4out_29_port, 
      PC_4out_28_port, PC_4out_27_port, PC_4out_26_port, PC_4out_25_port, 
      PC_4out_24_port, PC_4out_23_port, PC_4out_22_port, PC_4out_21_port, 
      PC_4out_20_port, PC_4out_19_port, PC_4out_18_port, PC_4out_17_port, 
      PC_4out_16_port, PC_4out_15_port, PC_4out_14_port, PC_4out_13_port, 
      PC_4out_12_port, PC_4out_11_port, PC_4out_10_port, PC_4out_9_port, 
      PC_4out_8_port, PC_4out_7_port, PC_4out_6_port, PC_4out_5_port, 
      PC_4out_4_port, PC_4out_3_port, PC_4out_2_port, PC_4out_1_port, 
      PC_4out_0_port );
   
   PC_REG : reg_N32_0 port map( clk => CLK, rst => RST, en => PC_EN, A(31) => 
                           IN_ID(31), A(30) => IN_ID(30), A(29) => IN_ID(29), 
                           A(28) => IN_ID(28), A(27) => IN_ID(27), A(26) => 
                           IN_ID(26), A(25) => IN_ID(25), A(24) => IN_ID(24), 
                           A(23) => IN_ID(23), A(22) => IN_ID(22), A(21) => 
                           IN_ID(21), A(20) => IN_ID(20), A(19) => IN_ID(19), 
                           A(18) => IN_ID(18), A(17) => IN_ID(17), A(16) => 
                           IN_ID(16), A(15) => IN_ID(15), A(14) => IN_ID(14), 
                           A(13) => IN_ID(13), A(12) => IN_ID(12), A(11) => 
                           IN_ID(11), A(10) => IN_ID(10), A(9) => IN_ID(9), 
                           A(8) => IN_ID(8), A(7) => IN_ID(7), A(6) => IN_ID(6)
                           , A(5) => IN_ID(5), A(4) => IN_ID(4), A(3) => 
                           IN_ID(3), A(2) => IN_ID(2), A(1) => IN_ID(1), A(0) 
                           => IN_ID(0), Y(31) => to_IRAM_31_port, Y(30) => 
                           to_IRAM_30_port, Y(29) => to_IRAM_29_port, Y(28) => 
                           to_IRAM_28_port, Y(27) => to_IRAM_27_port, Y(26) => 
                           to_IRAM_26_port, Y(25) => to_IRAM_25_port, Y(24) => 
                           to_IRAM_24_port, Y(23) => to_IRAM_23_port, Y(22) => 
                           to_IRAM_22_port, Y(21) => to_IRAM_21_port, Y(20) => 
                           to_IRAM_20_port, Y(19) => to_IRAM_19_port, Y(18) => 
                           to_IRAM_18_port, Y(17) => to_IRAM_17_port, Y(16) => 
                           to_IRAM_16_port, Y(15) => to_IRAM_15_port, Y(14) => 
                           to_IRAM_14_port, Y(13) => to_IRAM_13_port, Y(12) => 
                           to_IRAM_12_port, Y(11) => to_IRAM_11_port, Y(10) => 
                           to_IRAM_10_port, Y(9) => to_IRAM_9_port, Y(8) => 
                           to_IRAM_8_port, Y(7) => to_IRAM_7_port, Y(6) => 
                           to_IRAM_6_port, Y(5) => to_IRAM_5_port, Y(4) => 
                           to_IRAM_4_port, Y(3) => to_IRAM_3_port, Y(2) => 
                           to_IRAM_2_port, Y(1) => to_IRAM_1_port, Y(0) => 
                           to_IRAM_0_port);
   ADD : add4_NBIT32 port map( A(31) => to_IRAM_31_port, A(30) => 
                           to_IRAM_30_port, A(29) => to_IRAM_29_port, A(28) => 
                           to_IRAM_28_port, A(27) => to_IRAM_27_port, A(26) => 
                           to_IRAM_26_port, A(25) => to_IRAM_25_port, A(24) => 
                           to_IRAM_24_port, A(23) => to_IRAM_23_port, A(22) => 
                           to_IRAM_22_port, A(21) => to_IRAM_21_port, A(20) => 
                           to_IRAM_20_port, A(19) => to_IRAM_19_port, A(18) => 
                           to_IRAM_18_port, A(17) => to_IRAM_17_port, A(16) => 
                           to_IRAM_16_port, A(15) => to_IRAM_15_port, A(14) => 
                           to_IRAM_14_port, A(13) => to_IRAM_13_port, A(12) => 
                           to_IRAM_12_port, A(11) => to_IRAM_11_port, A(10) => 
                           to_IRAM_10_port, A(9) => to_IRAM_9_port, A(8) => 
                           to_IRAM_8_port, A(7) => to_IRAM_7_port, A(6) => 
                           to_IRAM_6_port, A(5) => to_IRAM_5_port, A(4) => 
                           to_IRAM_4_port, A(3) => to_IRAM_3_port, A(2) => 
                           to_IRAM_2_port, A(1) => to_IRAM_1_port, A(0) => 
                           to_IRAM_0_port, res(31) => PC_4out_31_port, res(30) 
                           => PC_4out_30_port, res(29) => PC_4out_29_port, 
                           res(28) => PC_4out_28_port, res(27) => 
                           PC_4out_27_port, res(26) => PC_4out_26_port, res(25)
                           => PC_4out_25_port, res(24) => PC_4out_24_port, 
                           res(23) => PC_4out_23_port, res(22) => 
                           PC_4out_22_port, res(21) => PC_4out_21_port, res(20)
                           => PC_4out_20_port, res(19) => PC_4out_19_port, 
                           res(18) => PC_4out_18_port, res(17) => 
                           PC_4out_17_port, res(16) => PC_4out_16_port, res(15)
                           => PC_4out_15_port, res(14) => PC_4out_14_port, 
                           res(13) => PC_4out_13_port, res(12) => 
                           PC_4out_12_port, res(11) => PC_4out_11_port, res(10)
                           => PC_4out_10_port, res(9) => PC_4out_9_port, res(8)
                           => PC_4out_8_port, res(7) => PC_4out_7_port, res(6) 
                           => PC_4out_6_port, res(5) => PC_4out_5_port, res(4) 
                           => PC_4out_4_port, res(3) => PC_4out_3_port, res(2) 
                           => PC_4out_2_port, res(1) => PC_4out_1_port, res(0) 
                           => PC_4out_0_port);
   NPC_REG : reg_N32_14 port map( clk => CLK, rst => RST, en => NPC_EN, A(31) 
                           => PC_4out_31_port, A(30) => PC_4out_30_port, A(29) 
                           => PC_4out_29_port, A(28) => PC_4out_28_port, A(27) 
                           => PC_4out_27_port, A(26) => PC_4out_26_port, A(25) 
                           => PC_4out_25_port, A(24) => PC_4out_24_port, A(23) 
                           => PC_4out_23_port, A(22) => PC_4out_22_port, A(21) 
                           => PC_4out_21_port, A(20) => PC_4out_20_port, A(19) 
                           => PC_4out_19_port, A(18) => PC_4out_18_port, A(17) 
                           => PC_4out_17_port, A(16) => PC_4out_16_port, A(15) 
                           => PC_4out_15_port, A(14) => PC_4out_14_port, A(13) 
                           => PC_4out_13_port, A(12) => PC_4out_12_port, A(11) 
                           => PC_4out_11_port, A(10) => PC_4out_10_port, A(9) 
                           => PC_4out_9_port, A(8) => PC_4out_8_port, A(7) => 
                           PC_4out_7_port, A(6) => PC_4out_6_port, A(5) => 
                           PC_4out_5_port, A(4) => PC_4out_4_port, A(3) => 
                           PC_4out_3_port, A(2) => PC_4out_2_port, A(1) => 
                           PC_4out_1_port, A(0) => PC_4out_0_port, Y(31) => 
                           NPC_out(31), Y(30) => NPC_out(30), Y(29) => 
                           NPC_out(29), Y(28) => NPC_out(28), Y(27) => 
                           NPC_out(27), Y(26) => NPC_out(26), Y(25) => 
                           NPC_out(25), Y(24) => NPC_out(24), Y(23) => 
                           NPC_out(23), Y(22) => NPC_out(22), Y(21) => 
                           NPC_out(21), Y(20) => NPC_out(20), Y(19) => 
                           NPC_out(19), Y(18) => NPC_out(18), Y(17) => 
                           NPC_out(17), Y(16) => NPC_out(16), Y(15) => 
                           NPC_out(15), Y(14) => NPC_out(14), Y(13) => 
                           NPC_out(13), Y(12) => NPC_out(12), Y(11) => 
                           NPC_out(11), Y(10) => NPC_out(10), Y(9) => 
                           NPC_out(9), Y(8) => NPC_out(8), Y(7) => NPC_out(7), 
                           Y(6) => NPC_out(6), Y(5) => NPC_out(5), Y(4) => 
                           NPC_out(4), Y(3) => NPC_out(3), Y(2) => NPC_out(2), 
                           Y(1) => NPC_out(1), Y(0) => NPC_out(0));
   I_REG : reg_N32_13 port map( clk => CLK, rst => RST, en => IR_EN, A(31) => 
                           from_IRAM(31), A(30) => from_IRAM(30), A(29) => 
                           from_IRAM(29), A(28) => from_IRAM(28), A(27) => 
                           from_IRAM(27), A(26) => from_IRAM(26), A(25) => 
                           from_IRAM(25), A(24) => from_IRAM(24), A(23) => 
                           from_IRAM(23), A(22) => from_IRAM(22), A(21) => 
                           from_IRAM(21), A(20) => from_IRAM(20), A(19) => 
                           from_IRAM(19), A(18) => from_IRAM(18), A(17) => 
                           from_IRAM(17), A(16) => from_IRAM(16), A(15) => 
                           from_IRAM(15), A(14) => from_IRAM(14), A(13) => 
                           from_IRAM(13), A(12) => from_IRAM(12), A(11) => 
                           from_IRAM(11), A(10) => from_IRAM(10), A(9) => 
                           from_IRAM(9), A(8) => from_IRAM(8), A(7) => 
                           from_IRAM(7), A(6) => from_IRAM(6), A(5) => 
                           from_IRAM(5), A(4) => from_IRAM(4), A(3) => 
                           from_IRAM(3), A(2) => from_IRAM(2), A(1) => 
                           from_IRAM(1), A(0) => from_IRAM(0), Y(31) => 
                           IREG_out(31), Y(30) => IREG_out(30), Y(29) => 
                           IREG_out(29), Y(28) => IREG_out(28), Y(27) => 
                           IREG_out(27), Y(26) => IREG_out(26), Y(25) => 
                           IREG_out(25), Y(24) => IREG_out(24), Y(23) => 
                           IREG_out(23), Y(22) => IREG_out(22), Y(21) => 
                           IREG_out(21), Y(20) => IREG_out(20), Y(19) => 
                           IREG_out(19), Y(18) => IREG_out(18), Y(17) => 
                           IREG_out(17), Y(16) => IREG_out(16), Y(15) => 
                           IREG_out(15), Y(14) => IREG_out(14), Y(13) => 
                           IREG_out(13), Y(12) => IREG_out(12), Y(11) => 
                           IREG_out(11), Y(10) => IREG_out(10), Y(9) => 
                           IREG_out(9), Y(8) => IREG_out(8), Y(7) => 
                           IREG_out(7), Y(6) => IREG_out(6), Y(5) => 
                           IREG_out(5), Y(4) => IREG_out(4), Y(3) => 
                           IREG_out(3), Y(2) => IREG_out(2), Y(1) => 
                           IREG_out(1), Y(0) => IREG_out(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE33_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE19 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         branch_taken : in std_logic;  IR_EN, NPC_EN, RegA_EN, RegB_EN, 
         RegIMM_EN, RT_REG_EN, IS_R_TYPE, J_EN, MUXA_SEL, MUXB_SEL, 
         ALU_OUTREG_EN, BRANCH_EN, BEQZ_OR_BNEZ, SH2_EN : out std_logic;  
         ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, LMD_EN, 
         WB_MUX_SEL, RF_WE, JAL_EN, PC_EN : out std_logic);

end dlx_cu_MICROCODE_MEM_SIZE33_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE19;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE33_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE19 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFR_X2
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic1_port, cw_FU_DU_10_port, cw_FU_DU_9_port, cw_FU_DU_8_port, 
      cw_FU_DU_7_port, cw_FU_DU_6_port, cw_FU_DU_5_port, cw_FU_DU_4_port, 
      cw_FU_DU_3_port, cw_FU_DU_2_port, cw_FU_DU_1_port, cw_FU_DU_0_port, 
      cw_EXU_4_port, cw_EXU_3_port, cw_EXU_2_port, cw_EXU_1_port, cw_EXU_0_port
      , cw_M_2_port, cw_M_1_port, cw_M_0_port, aluOpcode1_3_port, 
      aluOpcode1_2_port, aluOpcode1_1_port, aluOpcode1_0_port, N38, N39, N44, 
      N52, N56, N57, n411, n542, n582, n624, n717, n720, n28, n30, n32, n33, 
      n35, n37, n38_port, n39_port, n40, n41, n42, n43, n45, n52_port, n64, 
      net418894, net418895, net418897, net418900, net418907, net418910, 
      net421315, net421378, net421385, net421433, net421436, net421437, 
      net421439, net421458, net423241, net423243, net428488, net428487, 
      net428489, net428491, net428500, net428615, net428638, net428776, 
      net428766, net428758, net428753, net428744, net428742, net428738, 
      net428722, net428720, net428682, net428681, net428680, net428676, 
      net428860, net421452, net428617, net421454, net429511, net429479, 
      net429476, net428732, net428721, net428664, n61, n29, net427438, 
      net421457, net421456, net421311, net418906, n68, n67, n60, n53, net428858
      , net428684, net421441, net429500, net429469, net428734, net428497, 
      net423250, net423244, net423238, net421444, net421442, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, 
      n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672 : 
      std_logic;

begin
   PC_EN <= X_Logic1_port;
   
   X_Logic1_port <= '1';
   cw_FU_DU_reg_18_inst : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN 
                           => n794, Q => IR_EN, QN => n_1628);
   cw_FU_DU_reg_17_inst : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN 
                           => n796, Q => NPC_EN, QN => n_1629);
   cw_FU_DU_reg_15_inst : DFFR_X1 port map( D => net421378, CK => Clk, RN => 
                           n794, Q => RegB_EN, QN => n_1630);
   cw_FU_DU_reg_12_inst : DFFR_X1 port map( D => net421378, CK => Clk, RN => 
                           n794, Q => IS_R_TYPE, QN => n_1631);
   cw_FU_DU_reg_9_inst : DFFR_X1 port map( D => net421378, CK => Clk, RN => 
                           n797, Q => cw_FU_DU_9_port, QN => n_1632);
   cw_EXU_reg_9_inst : DFFR_X1 port map( D => cw_FU_DU_9_port, CK => Clk, RN =>
                           n797, Q => MUXB_SEL, QN => n_1633);
   cw_EXU_reg_8_inst : DFFR_X1 port map( D => cw_FU_DU_8_port, CK => Clk, RN =>
                           n797, Q => ALU_OUTREG_EN, QN => n_1634);
   cw_EXU_reg_7_inst : DFFR_X1 port map( D => cw_FU_DU_7_port, CK => Clk, RN =>
                           n797, Q => BRANCH_EN, QN => n_1635);
   cw_EXU_reg_6_inst : DFFR_X1 port map( D => cw_FU_DU_6_port, CK => Clk, RN =>
                           n796, Q => BEQZ_OR_BNEZ, QN => n_1636);
   cw_EXU_reg_5_inst : DFFR_X1 port map( D => cw_FU_DU_5_port, CK => Clk, RN =>
                           n796, Q => SH2_EN, QN => n_1637);
   cw_EXU_reg_4_inst : DFFR_X1 port map( D => cw_FU_DU_4_port, CK => Clk, RN =>
                           n796, Q => cw_EXU_4_port, QN => n_1638);
   cw_EXU_reg_3_inst : DFFR_X1 port map( D => cw_FU_DU_3_port, CK => Clk, RN =>
                           n795, Q => cw_EXU_3_port, QN => n_1639);
   cw_EXU_reg_2_inst : DFFR_X1 port map( D => cw_FU_DU_2_port, CK => Clk, RN =>
                           n796, Q => cw_EXU_2_port, QN => n_1640);
   cw_EXU_reg_1_inst : DFFR_X1 port map( D => cw_FU_DU_1_port, CK => Clk, RN =>
                           n796, Q => cw_EXU_1_port, QN => n_1641);
   cw_EXU_reg_0_inst : DFFR_X1 port map( D => cw_FU_DU_0_port, CK => Clk, RN =>
                           n796, Q => cw_EXU_0_port, QN => n_1642);
   cw_M_reg_4_inst : DFFR_X1 port map( D => cw_EXU_4_port, CK => Clk, RN => 
                           n796, Q => DRAM_WE, QN => n_1643);
   cw_M_reg_3_inst : DFFR_X1 port map( D => cw_EXU_3_port, CK => Clk, RN => 
                           n795, Q => LMD_EN, QN => n_1644);
   cw_M_reg_2_inst : DFFR_X1 port map( D => cw_EXU_2_port, CK => Clk, RN => 
                           n795, Q => cw_M_2_port, QN => n_1645);
   cw_M_reg_1_inst : DFFR_X1 port map( D => cw_EXU_1_port, CK => Clk, RN => 
                           n795, Q => cw_M_1_port, QN => n_1646);
   cw_M_reg_0_inst : DFFR_X1 port map( D => cw_EXU_0_port, CK => Clk, RN => 
                           n795, Q => cw_M_0_port, QN => n_1647);
   cw_WB_reg_2_inst : DFFR_X1 port map( D => cw_M_2_port, CK => Clk, RN => n795
                           , Q => WB_MUX_SEL, QN => n_1648);
   cw_WB_reg_1_inst : DFFR_X1 port map( D => cw_M_1_port, CK => Clk, RN => n795
                           , Q => RF_WE, QN => n_1649);
   cw_WB_reg_0_inst : DFFR_X1 port map( D => cw_M_0_port, CK => Clk, RN => n795
                           , Q => JAL_EN, QN => n_1650);
   aluOpcode2_reg_3_inst : DFFS_X1 port map( D => aluOpcode1_3_port, CK => Clk,
                           SN => n797, Q => ALU_OPCODE(0), QN => n_1651);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => aluOpcode1_2_port, CK => Clk,
                           RN => n795, Q => ALU_OPCODE(1), QN => n_1652);
   aluOpcode2_reg_1_inst : DFFS_X1 port map( D => aluOpcode1_1_port, CK => Clk,
                           SN => n797, Q => ALU_OPCODE(2), QN => n_1653);
   aluOpcode2_reg_0_inst : DFFS_X1 port map( D => aluOpcode1_0_port, CK => Clk,
                           SN => n797, Q => ALU_OPCODE(3), QN => n_1654);
   cw_EXU_reg_10_inst : DFFR_X1 port map( D => cw_FU_DU_10_port, CK => Clk, RN 
                           => n794, Q => MUXA_SEL, QN => n_1655);
   cw_FU_DU_reg_5_inst : DFFR_X1 port map( D => n765, CK => Clk, RN => n794, Q 
                           => cw_FU_DU_5_port, QN => n_1656);
   cw_FU_DU_reg_0_inst : DFFR_X1 port map( D => N38, CK => Clk, RN => n796, Q 
                           => cw_FU_DU_0_port, QN => n_1657);
   cw_FU_DU_reg_2_inst : DFFR_X1 port map( D => n542, CK => Clk, RN => n796, Q 
                           => cw_FU_DU_2_port, QN => n_1658);
   aluOpcode1_reg_1_inst : DFFS_X1 port map( D => N56, CK => Clk, SN => n797, Q
                           => aluOpcode1_1_port, QN => n_1659);
   U80 : XOR2_X1 port map( A => net418894, B => IR_IN(0), Z => n39_port);
   U82 : NAND3_X1 port map( A1 => n783, A2 => n35, A3 => n41, ZN => N56);
   aluOpcode1_reg_3_inst : DFFS_X1 port map( D => n717, CK => Clk, SN => n802, 
                           Q => aluOpcode1_3_port, QN => n_1660);
   aluOpcode1_reg_0_inst : DFFS_X1 port map( D => n720, CK => Clk, SN => n797, 
                           Q => aluOpcode1_0_port, QN => n_1661);
   cw_FU_DU_reg_4_inst : DFFR_X1 port map( D => net421385, CK => Clk, RN => 
                           n794, Q => cw_FU_DU_4_port, QN => n_1662);
   cw_FU_DU_reg_3_inst : DFFR_X1 port map( D => net421385, CK => Clk, RN => 
                           n795, Q => cw_FU_DU_3_port, QN => n_1663);
   cw_FU_DU_reg_11_inst : SDFFR_X1 port map( D => n791, SI => n792, SE => 
                           net421441, CK => Clk, RN => n795, Q => net423243, QN
                           => net428491);
   cw_FU_DU_reg_16_inst : SDFFR_X2 port map( D => N52, SI => n784, SE => 
                           net421378, CK => Clk, RN => n797, Q => RegA_EN, QN 
                           => n_1664);
   cw_FU_DU_reg_10_inst : DFFR_X2 port map( D => n582, CK => Clk, RN => n794, Q
                           => cw_FU_DU_10_port, QN => n_1665);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => N57, CK => Clk, RN => n794, Q
                           => aluOpcode1_2_port, QN => n_1666);
   cw_FU_DU_reg_6_inst : DFFR_X1 port map( D => N44, CK => Clk, RN => n797, Q 
                           => cw_FU_DU_6_port, QN => n_1667);
   cw_FU_DU_reg_8_inst : DFFR_X1 port map( D => n624, CK => Clk, RN => n797, Q 
                           => cw_FU_DU_8_port, QN => n_1668);
   cw_FU_DU_reg_13_inst : DFFR_X2 port map( D => n411, CK => Clk, RN => n794, Q
                           => RT_REG_EN, QN => n_1669);
   cw_FU_DU_reg_1_inst : DFFR_X2 port map( D => N39, CK => Clk, RN => n796, Q 
                           => cw_FU_DU_1_port, QN => n_1670);
   cw_FU_DU_reg_7_inst : DFFR_X1 port map( D => n765, CK => Clk, RN => n794, Q 
                           => cw_FU_DU_7_port, QN => n_1671);
   cw_FU_DU_reg_14_inst : DFFR_X2 port map( D => N52, CK => Clk, RN => n794, Q 
                           => RegIMM_EN, QN => n_1672);
   U3 : CLKBUF_X1 port map( A => net421441, Z => n764);
   U4 : NAND4_X1 port map( A1 => net418900, A2 => n67, A3 => net421452, A4 => 
                           net421439, ZN => net421457);
   U5 : NOR2_X1 port map( A1 => net418906, A2 => n776, ZN => n60);
   U6 : INV_X1 port map( A => net428721, ZN => n776);
   U7 : NAND2_X1 port map( A1 => net428681, A2 => net428682, ZN => net428680);
   U8 : INV_X1 port map( A => net421433, ZN => net428682);
   U9 : NOR2_X1 port map( A1 => IR_IN(28), A2 => IR_IN(30), ZN => net428681);
   U10 : NAND2_X1 port map( A1 => net429469, A2 => net429500, ZN => n775);
   U11 : INV_X1 port map( A => net421452, ZN => net429500);
   U12 : INV_X1 port map( A => IR_IN(28), ZN => net421311);
   U13 : INV_X1 port map( A => IR_IN(30), ZN => net429469);
   U14 : OAI21_X1 port map( B1 => n786, B2 => n787, A => IR_IN(27), ZN => 
                           net428738);
   U15 : NOR2_X1 port map( A1 => IR_IN(29), A2 => n38_port, ZN => n786);
   U16 : NOR2_X1 port map( A1 => n33, A2 => net421458, ZN => n787);
   U17 : AOI21_X1 port map( B1 => net428721, B2 => IR_IN(5), A => n780, ZN => 
                           net428720);
   U18 : NOR2_X1 port map( A1 => n40, A2 => IR_IN(0), ZN => n780);
   U19 : INV_X1 port map( A => n52_port, ZN => net428722);
   U20 : INV_X1 port map( A => net428680, ZN => net428684);
   U21 : NAND2_X1 port map( A1 => net428753, A2 => IR_IN(30), ZN => n789);
   U22 : INV_X1 port map( A => n45, ZN => net428753);
   U23 : NAND2_X1 port map( A1 => net428664, A2 => n52_port, ZN => n61);
   U24 : NOR2_X1 port map( A1 => net428680, A2 => IR_IN(26), ZN => net428664);
   U25 : INV_X1 port map( A => IR_IN(31), ZN => net429476);
   U26 : AND2_X1 port map( A1 => net428734, A2 => IR_IN(27), ZN => net429479);
   U27 : INV_X1 port map( A => n775, ZN => net428734);
   U28 : NAND2_X1 port map( A1 => net429469, A2 => IR_IN(28), ZN => n38_port);
   U29 : OAI21_X1 port map( B1 => IR_IN(1), B2 => n779, A => n781, ZN => 
                           net428721);
   U30 : NAND2_X1 port map( A1 => n778, A2 => net418897, ZN => n781);
   U31 : AOI21_X1 port map( B1 => IR_IN(3), B2 => IR_IN(0), A => IR_IN(2), ZN 
                           => n779);
   U32 : INV_X1 port map( A => IR_IN(0), ZN => n778);
   U33 : XNOR2_X1 port map( A => IR_IN(27), B => IR_IN(26), ZN => n37);
   U34 : OAI211_X1 port map( C1 => net418900, C2 => net429469, A => n68, B => 
                           net421439, ZN => n32);
   U35 : AND2_X1 port map( A1 => IR_IN(28), A2 => IR_IN(30), ZN => net428676);
   U36 : NOR2_X1 port map( A1 => net421433, A2 => IR_IN(26), ZN => n785);
   U37 : NAND2_X1 port map( A1 => net428742, A2 => n789, ZN => n788);
   U38 : OAI21_X1 port map( B1 => net428720, B2 => net428722, A => net428684, 
                           ZN => net428758);
   U39 : INV_X1 port map( A => n61, ZN => n777);
   U40 : INV_X1 port map( A => n29, ZN => net428732);
   U41 : NAND2_X1 port map( A1 => net429476, A2 => net421315, ZN => net421433);
   U42 : NOR2_X1 port map( A1 => net421433, A2 => IR_IN(27), ZN => n782);
   U43 : NAND2_X1 port map( A1 => IR_IN(30), A2 => net421439, ZN => net428488);
   U44 : NAND2_X1 port map( A1 => net428500, A2 => n766, ZN => net428615);
   U45 : AND2_X1 port map( A1 => net428500, A2 => n766, ZN => n765);
   U46 : INV_X1 port map( A => net428744, ZN => n35);
   U47 : OAI21_X1 port map( B1 => IR_IN(5), B2 => net428732, A => net418907, ZN
                           => net428744);
   U48 : AND2_X1 port map( A1 => n782, A2 => net421454, ZN => n766);
   U49 : AND2_X1 port map( A1 => IR_IN(5), A2 => n777, ZN => n767);
   U50 : NAND2_X1 port map( A1 => net429476, A2 => IR_IN(29), ZN => n33);
   U51 : NAND2_X1 port map( A1 => net428676, A2 => n785, ZN => net418907);
   U52 : AND2_X1 port map( A1 => IR_IN(27), A2 => net428684, ZN => n768);
   U53 : BUF_X1 port map( A => net429511, Z => n773);
   U54 : AND2_X1 port map( A1 => net428776, A2 => n790, ZN => n769);
   U55 : CLKBUF_X1 port map( A => net423241, Z => n770);
   U56 : AND2_X1 port map( A1 => net428858, A2 => n771, ZN => net428489);
   U57 : AND2_X1 port map( A1 => net428738, A2 => n790, ZN => n771);
   U58 : CLKBUF_X1 port map( A => net428491, Z => n772);
   U59 : NOR4_X1 port map( A1 => branch_taken, A2 => n775, A3 => net423243, A4 
                           => net418900, ZN => net423250);
   U60 : AND2_X1 port map( A1 => net421444, A2 => n53, ZN => net428497);
   U61 : AND2_X1 port map( A1 => net428491, A2 => n774, ZN => net428858);
   U62 : NAND4_X1 port map( A1 => net423241, A2 => net421441, A3 => net421444, 
                           A4 => net428617, ZN => N52);
   U63 : OAI211_X1 port map( C1 => n60, C2 => n29, A => net428491, B => n774, 
                           ZN => n53);
   U64 : INV_X1 port map( A => branch_taken, ZN => n774);
   U65 : AND2_X1 port map( A1 => net428497, A2 => net421442, ZN => net423238);
   U66 : NAND2_X1 port map( A1 => net423238, A2 => n764, ZN => n411);
   U67 : NAND2_X1 port map( A1 => net428497, A2 => net428615, ZN => n542);
   U68 : OAI21_X1 port map( B1 => net428860, B2 => IR_IN(29), A => net428497, 
                           ZN => N39);
   U69 : NAND2_X1 port map( A1 => net423250, A2 => IR_IN(31), ZN => net421442);
   U70 : NAND2_X1 port map( A1 => net423244, A2 => net421442, ZN => n582);
   U71 : AND2_X1 port map( A1 => net421444, A2 => n53, ZN => net423244);
   U72 : INV_X1 port map( A => n53, ZN => net421378);
   U73 : NAND2_X1 port map( A1 => net429511, A2 => IR_IN(31), ZN => net423241);
   U74 : NAND2_X1 port map( A1 => net427438, A2 => net421456, ZN => net421444);
   U75 : MUX2_X1 port map( A => IR_IN(27), B => net429476, S => net421452, Z =>
                           net428742);
   U76 : NAND2_X1 port map( A1 => net428858, A2 => n768, ZN => net421441);
   U77 : AND2_X1 port map( A1 => net428858, A2 => net428738, ZN => net428776);
   U78 : NOR2_X1 port map( A1 => net423243, A2 => branch_taken, ZN => net427438
                           );
   U79 : NOR2_X1 port map( A1 => branch_taken, A2 => net423243, ZN => net428500
                           );
   U81 : INV_X1 port map( A => n767, ZN => net418906);
   U83 : OR2_X1 port map( A1 => net418897, A2 => net418906, ZN => net428487);
   U84 : NOR2_X1 port map( A1 => n39_port, A2 => net418906, ZN => net421436);
   U85 : AOI221_X1 port map( B1 => IR_IN(1), B2 => n29, C1 => n30, C2 => n767, 
                           A => net418910, ZN => n28);
   U86 : AOI221_X1 port map( B1 => n29, B2 => net418894, C1 => n42, C2 => n767,
                           A => n43, ZN => n41);
   U87 : NAND3_X1 port map( A1 => n32, A2 => net418907, A3 => net421457, ZN => 
                           net421456);
   U88 : NAND2_X1 port map( A1 => IR_IN(30), A2 => net421311, ZN => n67);
   U89 : AOI221_X1 port map( B1 => IR_IN(26), B2 => net421315, C1 => IR_IN(29),
                           C2 => IR_IN(27), A => net421311, ZN => n45);
   U90 : AOI21_X1 port map( B1 => net418900, B2 => net421311, A => IR_IN(26), 
                           ZN => n68);
   U91 : NAND2_X1 port map( A1 => IR_IN(26), A2 => net421311, ZN => net421452);
   U92 : INV_X1 port map( A => IR_IN(27), ZN => net418900);
   U93 : AND2_X1 port map( A1 => net427438, A2 => net429479, ZN => net429511);
   U94 : NOR3_X1 port map( A1 => n40, A2 => IR_IN(0), A3 => n61, ZN => n29);
   U95 : INV_X1 port map( A => n40, ZN => net421437);
   U96 : NAND2_X1 port map( A1 => net428500, A2 => n766, ZN => net428617);
   U97 : INV_X1 port map( A => n773, ZN => net428860);
   U98 : INV_X1 port map( A => n38_port, ZN => net421454);
   U99 : AND2_X1 port map( A1 => net428776, A2 => n790, ZN => n783);
   n784 <= '1';
   U101 : INV_X1 port map( A => net428758, ZN => net428766);
   U102 : INV_X1 port map( A => net428500, ZN => net428638);
   U103 : NOR2_X1 port map( A1 => net428766, A2 => n788, ZN => n790);
   U104 : INV_X1 port map( A => n772, ZN => J_EN);
   U105 : NAND3_X1 port map( A1 => n769, A2 => net428488, A3 => net428487, ZN 
                           => n717);
   U106 : BUF_X1 port map( A => n793, Z => n798);
   U107 : BUF_X1 port map( A => n798, Z => n797);
   U108 : BUF_X1 port map( A => n799, Z => n794);
   U109 : BUF_X1 port map( A => n798, Z => n796);
   U110 : BUF_X1 port map( A => n799, Z => n795);
   U111 : BUF_X1 port map( A => n793, Z => n799);
   U112 : OAI211_X1 port map( C1 => net418900, C2 => net418907, A => net428489,
                           B => n28, ZN => n720);
   U113 : INV_X1 port map( A => n32, ZN => net418910);
   U114 : AOI21_X1 port map( B1 => net418895, B2 => net418894, A => IR_IN(0), 
                           ZN => n30);
   U115 : NOR2_X1 port map( A1 => IR_IN(2), A2 => net418897, ZN => n42);
   U116 : NOR4_X1 port map( A1 => IR_IN(27), A2 => IR_IN(26), A3 => n38_port, 
                           A4 => n33, ZN => n43);
   U117 : NOR4_X1 port map( A1 => IR_IN(6), A2 => IR_IN(4), A3 => IR_IN(10), A4
                           => n64, ZN => n52_port);
   U118 : OR4_X1 port map( A1 => IR_IN(8), A2 => IR_IN(7), A3 => IR_IN(27), A4 
                           => IR_IN(9), ZN => n64);
   U119 : NAND2_X1 port map( A1 => IR_IN(2), A2 => net418897, ZN => n40);
   U120 : INV_X1 port map( A => IR_IN(1), ZN => net418894);
   U121 : INV_X1 port map( A => IR_IN(3), ZN => net418897);
   U122 : BUF_X1 port map( A => n802, Z => n793);
   U123 : INV_X1 port map( A => IR_IN(2), ZN => net418895);
   n791 <= '1';
   n792 <= '0';
   U126 : OR2_X1 port map( A1 => n582, A2 => n765, ZN => n624);
   U127 : INV_X1 port map( A => IR_IN(29), ZN => net421315);
   U128 : INV_X1 port map( A => Rst, ZN => n802);
   U129 : INV_X1 port map( A => IR_IN(26), ZN => net421458);
   U130 : INV_X1 port map( A => n770, ZN => net421385);
   U131 : NOR2_X1 port map( A1 => n37, A2 => n38_port, ZN => n800);
   U132 : INV_X1 port map( A => n33, ZN => net421439);
   U133 : AOI221_X1 port map( B1 => net421436, B2 => net421437, C1 => n800, C2 
                           => net421439, A => net428744, ZN => n801);
   U134 : NOR2_X1 port map( A1 => net428638, A2 => n801, ZN => N57);
   U135 : NOR2_X1 port map( A1 => net428860, A2 => net421433, ZN => N38);
   U136 : NOR2_X1 port map( A1 => IR_IN(26), A2 => net428615, ZN => N44);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DATAPATH_N32 is

   port( CLK, RST : in std_logic;  ALU_FUNC : in std_logic_vector (0 to 3);  
         from_IRAM, from_DRAM : in std_logic_vector (31 downto 0);  IR_EN, 
         NPC_EN, RegA_EN, RegB_EN, RegIMM_EN, RT_REG_EN, IS_R_TYPE, J_EN, 
         MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, BRANCH_EN, BEQZ_OR_BNEZ, SH2_EN, 
         LMD_EN, WB_MUX_SEL, RF_WE, JAL_EN, PC_EN : in std_logic;  branch_taken
         : out std_logic;  addr_to_DRAM, data_to_DRAM, to_IRAM, IR : out 
         std_logic_vector (31 downto 0));

end DATAPATH_N32;

architecture SYN_STRUCTURAL of DATAPATH_N32 is

   component WBU_N32
      port( ALU_OUT, LOAD, NPC_REG_in, RT_REG_in : in std_logic_vector (31 
            downto 0);  IS_JAL, ALUOUT_OR_LOAD : in std_logic;  RF_ADDR, 
            RF_DATA : out std_logic_vector (31 downto 0));
   end component;
   
   component MU_N32
      port( CLK, RST, LMD_EN : in std_logic;  ALU_RESULT, RT_REG_in, NPC_REG_in
            , LMD_LATCH_in : in std_logic_vector (31 downto 0);  LMD_LATCH_out,
            ALU_REG_out, RT_REG_out, NPC_REG_out : out std_logic_vector (31 
            downto 0));
   end component;
   
   component EXU_N32
      port( CLK, RST, MUXA_SEL, MUXB_SEL, ZERO_EN, ZERO_SEL, ALUOUT_EN, 
            SHIFT2_EN : in std_logic;  ALU_FUNC : in std_logic_vector (0 to 3);
            NPC_REG, A_REG, B_REG, RT_REG, IMM_REG, PC_4 : in std_logic_vector 
            (31 downto 0);  ZERO : out std_logic;  BRANC_ADDR, ALU_OUT, 
            RT_REG_OUT, NPC_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component DU_N32
      port( J_EN, WR_EN, A_EN, B_EN, IMM_EN, RT_EN, is_R_type, BR_EN, clk, rst 
            : in std_logic;  NPC_IN, IR, DATAIN, ADDR_IN, BTA_OR_NPC : in 
            std_logic_vector (31 downto 0);  A, B, IMM, RT_OUT, NPC_OUT, PC_NXT
            : out std_logic_vector (31 downto 0));
   end component;
   
   component FU_N32
      port( CLK, RST, PC_EN, NPC_EN, IR_EN : in std_logic;  IN_ID, from_IRAM : 
            in std_logic_vector (31 downto 0);  to_IRAM, IREG_out, NPC_out, 
            PC_4out : out std_logic_vector (31 downto 0));
   end component;
   
   signal branch_taken_port, addr_to_DRAM_31_port, addr_to_DRAM_30_port, 
      addr_to_DRAM_29_port, addr_to_DRAM_28_port, addr_to_DRAM_27_port, 
      addr_to_DRAM_26_port, addr_to_DRAM_25_port, addr_to_DRAM_24_port, 
      addr_to_DRAM_23_port, addr_to_DRAM_22_port, addr_to_DRAM_21_port, 
      addr_to_DRAM_20_port, addr_to_DRAM_19_port, addr_to_DRAM_18_port, 
      addr_to_DRAM_17_port, addr_to_DRAM_16_port, addr_to_DRAM_15_port, 
      addr_to_DRAM_14_port, addr_to_DRAM_13_port, addr_to_DRAM_12_port, 
      addr_to_DRAM_11_port, addr_to_DRAM_10_port, addr_to_DRAM_9_port, 
      addr_to_DRAM_8_port, addr_to_DRAM_7_port, addr_to_DRAM_6_port, 
      addr_to_DRAM_5_port, addr_to_DRAM_4_port, addr_to_DRAM_3_port, 
      addr_to_DRAM_2_port, addr_to_DRAM_1_port, addr_to_DRAM_0_port, 
      data_to_DRAM_31_port, data_to_DRAM_30_port, data_to_DRAM_29_port, 
      data_to_DRAM_28_port, data_to_DRAM_27_port, data_to_DRAM_26_port, 
      data_to_DRAM_25_port, data_to_DRAM_24_port, data_to_DRAM_23_port, 
      data_to_DRAM_22_port, data_to_DRAM_21_port, data_to_DRAM_20_port, 
      data_to_DRAM_19_port, data_to_DRAM_18_port, data_to_DRAM_17_port, 
      data_to_DRAM_16_port, data_to_DRAM_15_port, data_to_DRAM_14_port, 
      data_to_DRAM_13_port, data_to_DRAM_12_port, data_to_DRAM_11_port, 
      data_to_DRAM_10_port, data_to_DRAM_9_port, data_to_DRAM_8_port, 
      data_to_DRAM_7_port, data_to_DRAM_6_port, data_to_DRAM_5_port, 
      data_to_DRAM_4_port, data_to_DRAM_3_port, data_to_DRAM_2_port, 
      data_to_DRAM_1_port, data_to_DRAM_0_port, IR_31_port, IR_30_port, 
      IR_29_port, IR_28_port, IR_27_port, IR_26_port, IR_25_port, IR_24_port, 
      IR_23_port, IR_22_port, IR_21_port, IR_20_port, IR_19_port, IR_18_port, 
      IR_17_port, IR_16_port, IR_15_port, IR_14_port, IR_13_port, IR_12_port, 
      IR_11_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, IR_6_port, 
      IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, IR_0_port, 
      pc_nxt_s_31_port, pc_nxt_s_30_port, pc_nxt_s_29_port, pc_nxt_s_28_port, 
      pc_nxt_s_27_port, pc_nxt_s_26_port, pc_nxt_s_25_port, pc_nxt_s_24_port, 
      pc_nxt_s_23_port, pc_nxt_s_22_port, pc_nxt_s_21_port, pc_nxt_s_20_port, 
      pc_nxt_s_19_port, pc_nxt_s_18_port, pc_nxt_s_17_port, pc_nxt_s_16_port, 
      pc_nxt_s_15_port, pc_nxt_s_14_port, pc_nxt_s_13_port, pc_nxt_s_12_port, 
      pc_nxt_s_11_port, pc_nxt_s_10_port, pc_nxt_s_9_port, pc_nxt_s_8_port, 
      pc_nxt_s_7_port, pc_nxt_s_6_port, pc_nxt_s_5_port, pc_nxt_s_4_port, 
      pc_nxt_s_3_port, pc_nxt_s_2_port, pc_nxt_s_1_port, pc_nxt_s_0_port, 
      npc_reg1_s_31_port, npc_reg1_s_30_port, npc_reg1_s_29_port, 
      npc_reg1_s_28_port, npc_reg1_s_27_port, npc_reg1_s_26_port, 
      npc_reg1_s_25_port, npc_reg1_s_24_port, npc_reg1_s_23_port, 
      npc_reg1_s_22_port, npc_reg1_s_21_port, npc_reg1_s_20_port, 
      npc_reg1_s_19_port, npc_reg1_s_18_port, npc_reg1_s_17_port, 
      npc_reg1_s_16_port, npc_reg1_s_15_port, npc_reg1_s_14_port, 
      npc_reg1_s_13_port, npc_reg1_s_12_port, npc_reg1_s_11_port, 
      npc_reg1_s_10_port, npc_reg1_s_9_port, npc_reg1_s_8_port, 
      npc_reg1_s_7_port, npc_reg1_s_6_port, npc_reg1_s_5_port, 
      npc_reg1_s_4_port, npc_reg1_s_3_port, npc_reg1_s_2_port, 
      npc_reg1_s_1_port, npc_reg1_s_0_port, pc4_s_31_port, pc4_s_30_port, 
      pc4_s_29_port, pc4_s_28_port, pc4_s_27_port, pc4_s_26_port, pc4_s_25_port
      , pc4_s_24_port, pc4_s_23_port, pc4_s_22_port, pc4_s_21_port, 
      pc4_s_20_port, pc4_s_19_port, pc4_s_18_port, pc4_s_17_port, pc4_s_16_port
      , pc4_s_15_port, pc4_s_14_port, pc4_s_13_port, pc4_s_12_port, 
      pc4_s_11_port, pc4_s_10_port, pc4_s_9_port, pc4_s_8_port, pc4_s_7_port, 
      pc4_s_6_port, pc4_s_5_port, pc4_s_4_port, pc4_s_3_port, pc4_s_2_port, 
      pc4_s_1_port, pc4_s_0_port, wb_data_s_31_port, wb_data_s_30_port, 
      wb_data_s_29_port, wb_data_s_28_port, wb_data_s_27_port, 
      wb_data_s_26_port, wb_data_s_25_port, wb_data_s_24_port, 
      wb_data_s_23_port, wb_data_s_22_port, wb_data_s_21_port, 
      wb_data_s_20_port, wb_data_s_19_port, wb_data_s_18_port, 
      wb_data_s_17_port, wb_data_s_16_port, wb_data_s_15_port, 
      wb_data_s_14_port, wb_data_s_13_port, wb_data_s_12_port, 
      wb_data_s_11_port, wb_data_s_10_port, wb_data_s_9_port, wb_data_s_8_port,
      wb_data_s_7_port, wb_data_s_6_port, wb_data_s_5_port, wb_data_s_4_port, 
      wb_data_s_3_port, wb_data_s_2_port, wb_data_s_1_port, wb_data_s_0_port, 
      wb_addr_s_31_port, wb_addr_s_30_port, wb_addr_s_29_port, 
      wb_addr_s_28_port, wb_addr_s_27_port, wb_addr_s_26_port, 
      wb_addr_s_25_port, wb_addr_s_24_port, wb_addr_s_23_port, 
      wb_addr_s_22_port, wb_addr_s_21_port, wb_addr_s_20_port, 
      wb_addr_s_19_port, wb_addr_s_18_port, wb_addr_s_17_port, 
      wb_addr_s_16_port, wb_addr_s_15_port, wb_addr_s_14_port, 
      wb_addr_s_13_port, wb_addr_s_12_port, wb_addr_s_11_port, 
      wb_addr_s_10_port, wb_addr_s_9_port, wb_addr_s_8_port, wb_addr_s_7_port, 
      wb_addr_s_6_port, wb_addr_s_5_port, wb_addr_s_4_port, wb_addr_s_3_port, 
      wb_addr_s_2_port, wb_addr_s_1_port, wb_addr_s_0_port, b_addr_s_31_port, 
      b_addr_s_30_port, b_addr_s_29_port, b_addr_s_28_port, b_addr_s_27_port, 
      b_addr_s_26_port, b_addr_s_25_port, b_addr_s_24_port, b_addr_s_23_port, 
      b_addr_s_22_port, b_addr_s_21_port, b_addr_s_20_port, b_addr_s_19_port, 
      b_addr_s_18_port, b_addr_s_17_port, b_addr_s_16_port, b_addr_s_15_port, 
      b_addr_s_14_port, b_addr_s_13_port, b_addr_s_12_port, b_addr_s_11_port, 
      b_addr_s_10_port, b_addr_s_9_port, b_addr_s_8_port, b_addr_s_7_port, 
      b_addr_s_6_port, b_addr_s_5_port, b_addr_s_4_port, b_addr_s_3_port, 
      b_addr_s_2_port, b_addr_s_1_port, b_addr_s_0_port, a_reg_s_31_port, 
      a_reg_s_30_port, a_reg_s_29_port, a_reg_s_28_port, a_reg_s_27_port, 
      a_reg_s_26_port, a_reg_s_25_port, a_reg_s_24_port, a_reg_s_23_port, 
      a_reg_s_22_port, a_reg_s_21_port, a_reg_s_20_port, a_reg_s_19_port, 
      a_reg_s_18_port, a_reg_s_17_port, a_reg_s_16_port, a_reg_s_15_port, 
      a_reg_s_14_port, a_reg_s_13_port, a_reg_s_12_port, a_reg_s_11_port, 
      a_reg_s_10_port, a_reg_s_9_port, a_reg_s_8_port, a_reg_s_7_port, 
      a_reg_s_6_port, a_reg_s_5_port, a_reg_s_4_port, a_reg_s_3_port, 
      a_reg_s_2_port, a_reg_s_1_port, a_reg_s_0_port, b_reg_s_31_port, 
      b_reg_s_30_port, b_reg_s_29_port, b_reg_s_28_port, b_reg_s_27_port, 
      b_reg_s_26_port, b_reg_s_25_port, b_reg_s_24_port, b_reg_s_23_port, 
      b_reg_s_22_port, b_reg_s_21_port, b_reg_s_20_port, b_reg_s_19_port, 
      b_reg_s_18_port, b_reg_s_17_port, b_reg_s_16_port, b_reg_s_15_port, 
      b_reg_s_14_port, b_reg_s_13_port, b_reg_s_12_port, b_reg_s_11_port, 
      b_reg_s_10_port, b_reg_s_9_port, b_reg_s_8_port, b_reg_s_7_port, 
      b_reg_s_6_port, b_reg_s_5_port, b_reg_s_4_port, b_reg_s_3_port, 
      b_reg_s_2_port, b_reg_s_1_port, b_reg_s_0_port, imm_reg_s_31_port, 
      imm_reg_s_30_port, imm_reg_s_29_port, imm_reg_s_28_port, 
      imm_reg_s_27_port, imm_reg_s_26_port, imm_reg_s_25_port, 
      imm_reg_s_24_port, imm_reg_s_23_port, imm_reg_s_22_port, 
      imm_reg_s_21_port, imm_reg_s_20_port, imm_reg_s_19_port, 
      imm_reg_s_18_port, imm_reg_s_17_port, imm_reg_s_16_port, 
      imm_reg_s_15_port, imm_reg_s_14_port, imm_reg_s_13_port, 
      imm_reg_s_12_port, imm_reg_s_11_port, imm_reg_s_10_port, imm_reg_s_9_port
      , imm_reg_s_8_port, imm_reg_s_7_port, imm_reg_s_6_port, imm_reg_s_5_port,
      imm_reg_s_4_port, imm_reg_s_3_port, imm_reg_s_2_port, imm_reg_s_1_port, 
      imm_reg_s_0_port, rt_reg1_s_31_port, rt_reg1_s_30_port, rt_reg1_s_29_port
      , rt_reg1_s_28_port, rt_reg1_s_27_port, rt_reg1_s_26_port, 
      rt_reg1_s_25_port, rt_reg1_s_24_port, rt_reg1_s_23_port, 
      rt_reg1_s_22_port, rt_reg1_s_21_port, rt_reg1_s_20_port, 
      rt_reg1_s_19_port, rt_reg1_s_18_port, rt_reg1_s_17_port, 
      rt_reg1_s_16_port, rt_reg1_s_15_port, rt_reg1_s_14_port, 
      rt_reg1_s_13_port, rt_reg1_s_12_port, rt_reg1_s_11_port, 
      rt_reg1_s_10_port, rt_reg1_s_9_port, rt_reg1_s_8_port, rt_reg1_s_7_port, 
      rt_reg1_s_6_port, rt_reg1_s_5_port, rt_reg1_s_4_port, rt_reg1_s_3_port, 
      rt_reg1_s_2_port, rt_reg1_s_1_port, rt_reg1_s_0_port, npc_reg2_s_31_port,
      npc_reg2_s_30_port, npc_reg2_s_29_port, npc_reg2_s_28_port, 
      npc_reg2_s_27_port, npc_reg2_s_26_port, npc_reg2_s_25_port, 
      npc_reg2_s_24_port, npc_reg2_s_23_port, npc_reg2_s_22_port, 
      npc_reg2_s_21_port, npc_reg2_s_20_port, npc_reg2_s_19_port, 
      npc_reg2_s_18_port, npc_reg2_s_17_port, npc_reg2_s_16_port, 
      npc_reg2_s_15_port, npc_reg2_s_14_port, npc_reg2_s_13_port, 
      npc_reg2_s_12_port, npc_reg2_s_11_port, npc_reg2_s_10_port, 
      npc_reg2_s_9_port, npc_reg2_s_8_port, npc_reg2_s_7_port, 
      npc_reg2_s_6_port, npc_reg2_s_5_port, npc_reg2_s_4_port, 
      npc_reg2_s_3_port, npc_reg2_s_2_port, npc_reg2_s_1_port, 
      npc_reg2_s_0_port, npc_reg3_s_31_port, npc_reg3_s_30_port, 
      npc_reg3_s_29_port, npc_reg3_s_28_port, npc_reg3_s_27_port, 
      npc_reg3_s_26_port, npc_reg3_s_25_port, npc_reg3_s_24_port, 
      npc_reg3_s_23_port, npc_reg3_s_22_port, npc_reg3_s_21_port, 
      npc_reg3_s_20_port, npc_reg3_s_19_port, npc_reg3_s_18_port, 
      npc_reg3_s_17_port, npc_reg3_s_16_port, npc_reg3_s_15_port, 
      npc_reg3_s_14_port, npc_reg3_s_13_port, npc_reg3_s_12_port, 
      npc_reg3_s_11_port, npc_reg3_s_10_port, npc_reg3_s_9_port, 
      npc_reg3_s_8_port, npc_reg3_s_7_port, npc_reg3_s_6_port, 
      npc_reg3_s_5_port, npc_reg3_s_4_port, npc_reg3_s_3_port, 
      npc_reg3_s_2_port, npc_reg3_s_1_port, npc_reg3_s_0_port, 
      lmd_out_s_31_port, lmd_out_s_30_port, lmd_out_s_29_port, 
      lmd_out_s_28_port, lmd_out_s_27_port, lmd_out_s_26_port, 
      lmd_out_s_25_port, lmd_out_s_24_port, lmd_out_s_23_port, 
      lmd_out_s_22_port, lmd_out_s_21_port, lmd_out_s_20_port, 
      lmd_out_s_19_port, lmd_out_s_18_port, lmd_out_s_17_port, 
      lmd_out_s_16_port, lmd_out_s_15_port, lmd_out_s_14_port, 
      lmd_out_s_13_port, lmd_out_s_12_port, lmd_out_s_11_port, 
      lmd_out_s_10_port, lmd_out_s_9_port, lmd_out_s_8_port, lmd_out_s_7_port, 
      lmd_out_s_6_port, lmd_out_s_5_port, lmd_out_s_4_port, lmd_out_s_3_port, 
      lmd_out_s_2_port, lmd_out_s_1_port, lmd_out_s_0_port, alu_out2_s_31_port,
      alu_out2_s_30_port, alu_out2_s_29_port, alu_out2_s_28_port, 
      alu_out2_s_27_port, alu_out2_s_26_port, alu_out2_s_25_port, 
      alu_out2_s_24_port, alu_out2_s_23_port, alu_out2_s_22_port, 
      alu_out2_s_21_port, alu_out2_s_20_port, alu_out2_s_19_port, 
      alu_out2_s_18_port, alu_out2_s_17_port, alu_out2_s_16_port, 
      alu_out2_s_15_port, alu_out2_s_14_port, alu_out2_s_13_port, 
      alu_out2_s_12_port, alu_out2_s_11_port, alu_out2_s_10_port, 
      alu_out2_s_9_port, alu_out2_s_8_port, alu_out2_s_7_port, 
      alu_out2_s_6_port, alu_out2_s_5_port, alu_out2_s_4_port, 
      alu_out2_s_3_port, alu_out2_s_2_port, alu_out2_s_1_port, 
      alu_out2_s_0_port, rt_reg3_s_31_port, rt_reg3_s_30_port, 
      rt_reg3_s_29_port, rt_reg3_s_28_port, rt_reg3_s_27_port, 
      rt_reg3_s_26_port, rt_reg3_s_25_port, rt_reg3_s_24_port, 
      rt_reg3_s_23_port, rt_reg3_s_22_port, rt_reg3_s_21_port, 
      rt_reg3_s_20_port, rt_reg3_s_19_port, rt_reg3_s_18_port, 
      rt_reg3_s_17_port, rt_reg3_s_16_port, rt_reg3_s_15_port, 
      rt_reg3_s_14_port, rt_reg3_s_13_port, rt_reg3_s_12_port, 
      rt_reg3_s_11_port, rt_reg3_s_10_port, rt_reg3_s_9_port, rt_reg3_s_8_port,
      rt_reg3_s_7_port, rt_reg3_s_6_port, rt_reg3_s_5_port, rt_reg3_s_4_port, 
      rt_reg3_s_3_port, rt_reg3_s_2_port, rt_reg3_s_1_port, rt_reg3_s_0_port, 
      npc_reg4_s_31_port, npc_reg4_s_30_port, npc_reg4_s_29_port, 
      npc_reg4_s_28_port, npc_reg4_s_27_port, npc_reg4_s_26_port, 
      npc_reg4_s_25_port, npc_reg4_s_24_port, npc_reg4_s_23_port, 
      npc_reg4_s_22_port, npc_reg4_s_21_port, npc_reg4_s_20_port, 
      npc_reg4_s_19_port, npc_reg4_s_18_port, npc_reg4_s_17_port, 
      npc_reg4_s_16_port, npc_reg4_s_15_port, npc_reg4_s_14_port, 
      npc_reg4_s_13_port, npc_reg4_s_12_port, npc_reg4_s_11_port, 
      npc_reg4_s_10_port, npc_reg4_s_9_port, npc_reg4_s_8_port, 
      npc_reg4_s_7_port, npc_reg4_s_6_port, npc_reg4_s_5_port, 
      npc_reg4_s_4_port, npc_reg4_s_3_port, npc_reg4_s_2_port, 
      npc_reg4_s_1_port, npc_reg4_s_0_port : std_logic;

begin
   branch_taken <= branch_taken_port;
   addr_to_DRAM <= ( addr_to_DRAM_31_port, addr_to_DRAM_30_port, 
      addr_to_DRAM_29_port, addr_to_DRAM_28_port, addr_to_DRAM_27_port, 
      addr_to_DRAM_26_port, addr_to_DRAM_25_port, addr_to_DRAM_24_port, 
      addr_to_DRAM_23_port, addr_to_DRAM_22_port, addr_to_DRAM_21_port, 
      addr_to_DRAM_20_port, addr_to_DRAM_19_port, addr_to_DRAM_18_port, 
      addr_to_DRAM_17_port, addr_to_DRAM_16_port, addr_to_DRAM_15_port, 
      addr_to_DRAM_14_port, addr_to_DRAM_13_port, addr_to_DRAM_12_port, 
      addr_to_DRAM_11_port, addr_to_DRAM_10_port, addr_to_DRAM_9_port, 
      addr_to_DRAM_8_port, addr_to_DRAM_7_port, addr_to_DRAM_6_port, 
      addr_to_DRAM_5_port, addr_to_DRAM_4_port, addr_to_DRAM_3_port, 
      addr_to_DRAM_2_port, addr_to_DRAM_1_port, addr_to_DRAM_0_port );
   data_to_DRAM <= ( data_to_DRAM_31_port, data_to_DRAM_30_port, 
      data_to_DRAM_29_port, data_to_DRAM_28_port, data_to_DRAM_27_port, 
      data_to_DRAM_26_port, data_to_DRAM_25_port, data_to_DRAM_24_port, 
      data_to_DRAM_23_port, data_to_DRAM_22_port, data_to_DRAM_21_port, 
      data_to_DRAM_20_port, data_to_DRAM_19_port, data_to_DRAM_18_port, 
      data_to_DRAM_17_port, data_to_DRAM_16_port, data_to_DRAM_15_port, 
      data_to_DRAM_14_port, data_to_DRAM_13_port, data_to_DRAM_12_port, 
      data_to_DRAM_11_port, data_to_DRAM_10_port, data_to_DRAM_9_port, 
      data_to_DRAM_8_port, data_to_DRAM_7_port, data_to_DRAM_6_port, 
      data_to_DRAM_5_port, data_to_DRAM_4_port, data_to_DRAM_3_port, 
      data_to_DRAM_2_port, data_to_DRAM_1_port, data_to_DRAM_0_port );
   IR <= ( IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, 
      IR_20_port, IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, 
      IR_14_port, IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, 
      IR_8_port, IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, 
      IR_2_port, IR_1_port, IR_0_port );
   
   F_STAGE : FU_N32 port map( CLK => CLK, RST => RST, PC_EN => PC_EN, NPC_EN =>
                           NPC_EN, IR_EN => IR_EN, IN_ID(31) => 
                           pc_nxt_s_31_port, IN_ID(30) => pc_nxt_s_30_port, 
                           IN_ID(29) => pc_nxt_s_29_port, IN_ID(28) => 
                           pc_nxt_s_28_port, IN_ID(27) => pc_nxt_s_27_port, 
                           IN_ID(26) => pc_nxt_s_26_port, IN_ID(25) => 
                           pc_nxt_s_25_port, IN_ID(24) => pc_nxt_s_24_port, 
                           IN_ID(23) => pc_nxt_s_23_port, IN_ID(22) => 
                           pc_nxt_s_22_port, IN_ID(21) => pc_nxt_s_21_port, 
                           IN_ID(20) => pc_nxt_s_20_port, IN_ID(19) => 
                           pc_nxt_s_19_port, IN_ID(18) => pc_nxt_s_18_port, 
                           IN_ID(17) => pc_nxt_s_17_port, IN_ID(16) => 
                           pc_nxt_s_16_port, IN_ID(15) => pc_nxt_s_15_port, 
                           IN_ID(14) => pc_nxt_s_14_port, IN_ID(13) => 
                           pc_nxt_s_13_port, IN_ID(12) => pc_nxt_s_12_port, 
                           IN_ID(11) => pc_nxt_s_11_port, IN_ID(10) => 
                           pc_nxt_s_10_port, IN_ID(9) => pc_nxt_s_9_port, 
                           IN_ID(8) => pc_nxt_s_8_port, IN_ID(7) => 
                           pc_nxt_s_7_port, IN_ID(6) => pc_nxt_s_6_port, 
                           IN_ID(5) => pc_nxt_s_5_port, IN_ID(4) => 
                           pc_nxt_s_4_port, IN_ID(3) => pc_nxt_s_3_port, 
                           IN_ID(2) => pc_nxt_s_2_port, IN_ID(1) => 
                           pc_nxt_s_1_port, IN_ID(0) => pc_nxt_s_0_port, 
                           from_IRAM(31) => from_IRAM(31), from_IRAM(30) => 
                           from_IRAM(30), from_IRAM(29) => from_IRAM(29), 
                           from_IRAM(28) => from_IRAM(28), from_IRAM(27) => 
                           from_IRAM(27), from_IRAM(26) => from_IRAM(26), 
                           from_IRAM(25) => from_IRAM(25), from_IRAM(24) => 
                           from_IRAM(24), from_IRAM(23) => from_IRAM(23), 
                           from_IRAM(22) => from_IRAM(22), from_IRAM(21) => 
                           from_IRAM(21), from_IRAM(20) => from_IRAM(20), 
                           from_IRAM(19) => from_IRAM(19), from_IRAM(18) => 
                           from_IRAM(18), from_IRAM(17) => from_IRAM(17), 
                           from_IRAM(16) => from_IRAM(16), from_IRAM(15) => 
                           from_IRAM(15), from_IRAM(14) => from_IRAM(14), 
                           from_IRAM(13) => from_IRAM(13), from_IRAM(12) => 
                           from_IRAM(12), from_IRAM(11) => from_IRAM(11), 
                           from_IRAM(10) => from_IRAM(10), from_IRAM(9) => 
                           from_IRAM(9), from_IRAM(8) => from_IRAM(8), 
                           from_IRAM(7) => from_IRAM(7), from_IRAM(6) => 
                           from_IRAM(6), from_IRAM(5) => from_IRAM(5), 
                           from_IRAM(4) => from_IRAM(4), from_IRAM(3) => 
                           from_IRAM(3), from_IRAM(2) => from_IRAM(2), 
                           from_IRAM(1) => from_IRAM(1), from_IRAM(0) => 
                           from_IRAM(0), to_IRAM(31) => to_IRAM(31), 
                           to_IRAM(30) => to_IRAM(30), to_IRAM(29) => 
                           to_IRAM(29), to_IRAM(28) => to_IRAM(28), to_IRAM(27)
                           => to_IRAM(27), to_IRAM(26) => to_IRAM(26), 
                           to_IRAM(25) => to_IRAM(25), to_IRAM(24) => 
                           to_IRAM(24), to_IRAM(23) => to_IRAM(23), to_IRAM(22)
                           => to_IRAM(22), to_IRAM(21) => to_IRAM(21), 
                           to_IRAM(20) => to_IRAM(20), to_IRAM(19) => 
                           to_IRAM(19), to_IRAM(18) => to_IRAM(18), to_IRAM(17)
                           => to_IRAM(17), to_IRAM(16) => to_IRAM(16), 
                           to_IRAM(15) => to_IRAM(15), to_IRAM(14) => 
                           to_IRAM(14), to_IRAM(13) => to_IRAM(13), to_IRAM(12)
                           => to_IRAM(12), to_IRAM(11) => to_IRAM(11), 
                           to_IRAM(10) => to_IRAM(10), to_IRAM(9) => to_IRAM(9)
                           , to_IRAM(8) => to_IRAM(8), to_IRAM(7) => to_IRAM(7)
                           , to_IRAM(6) => to_IRAM(6), to_IRAM(5) => to_IRAM(5)
                           , to_IRAM(4) => to_IRAM(4), to_IRAM(3) => to_IRAM(3)
                           , to_IRAM(2) => to_IRAM(2), to_IRAM(1) => to_IRAM(1)
                           , to_IRAM(0) => to_IRAM(0), IREG_out(31) => 
                           IR_31_port, IREG_out(30) => IR_30_port, IREG_out(29)
                           => IR_29_port, IREG_out(28) => IR_28_port, 
                           IREG_out(27) => IR_27_port, IREG_out(26) => 
                           IR_26_port, IREG_out(25) => IR_25_port, IREG_out(24)
                           => IR_24_port, IREG_out(23) => IR_23_port, 
                           IREG_out(22) => IR_22_port, IREG_out(21) => 
                           IR_21_port, IREG_out(20) => IR_20_port, IREG_out(19)
                           => IR_19_port, IREG_out(18) => IR_18_port, 
                           IREG_out(17) => IR_17_port, IREG_out(16) => 
                           IR_16_port, IREG_out(15) => IR_15_port, IREG_out(14)
                           => IR_14_port, IREG_out(13) => IR_13_port, 
                           IREG_out(12) => IR_12_port, IREG_out(11) => 
                           IR_11_port, IREG_out(10) => IR_10_port, IREG_out(9) 
                           => IR_9_port, IREG_out(8) => IR_8_port, IREG_out(7) 
                           => IR_7_port, IREG_out(6) => IR_6_port, IREG_out(5) 
                           => IR_5_port, IREG_out(4) => IR_4_port, IREG_out(3) 
                           => IR_3_port, IREG_out(2) => IR_2_port, IREG_out(1) 
                           => IR_1_port, IREG_out(0) => IR_0_port, NPC_out(31) 
                           => npc_reg1_s_31_port, NPC_out(30) => 
                           npc_reg1_s_30_port, NPC_out(29) => 
                           npc_reg1_s_29_port, NPC_out(28) => 
                           npc_reg1_s_28_port, NPC_out(27) => 
                           npc_reg1_s_27_port, NPC_out(26) => 
                           npc_reg1_s_26_port, NPC_out(25) => 
                           npc_reg1_s_25_port, NPC_out(24) => 
                           npc_reg1_s_24_port, NPC_out(23) => 
                           npc_reg1_s_23_port, NPC_out(22) => 
                           npc_reg1_s_22_port, NPC_out(21) => 
                           npc_reg1_s_21_port, NPC_out(20) => 
                           npc_reg1_s_20_port, NPC_out(19) => 
                           npc_reg1_s_19_port, NPC_out(18) => 
                           npc_reg1_s_18_port, NPC_out(17) => 
                           npc_reg1_s_17_port, NPC_out(16) => 
                           npc_reg1_s_16_port, NPC_out(15) => 
                           npc_reg1_s_15_port, NPC_out(14) => 
                           npc_reg1_s_14_port, NPC_out(13) => 
                           npc_reg1_s_13_port, NPC_out(12) => 
                           npc_reg1_s_12_port, NPC_out(11) => 
                           npc_reg1_s_11_port, NPC_out(10) => 
                           npc_reg1_s_10_port, NPC_out(9) => npc_reg1_s_9_port,
                           NPC_out(8) => npc_reg1_s_8_port, NPC_out(7) => 
                           npc_reg1_s_7_port, NPC_out(6) => npc_reg1_s_6_port, 
                           NPC_out(5) => npc_reg1_s_5_port, NPC_out(4) => 
                           npc_reg1_s_4_port, NPC_out(3) => npc_reg1_s_3_port, 
                           NPC_out(2) => npc_reg1_s_2_port, NPC_out(1) => 
                           npc_reg1_s_1_port, NPC_out(0) => npc_reg1_s_0_port, 
                           PC_4out(31) => pc4_s_31_port, PC_4out(30) => 
                           pc4_s_30_port, PC_4out(29) => pc4_s_29_port, 
                           PC_4out(28) => pc4_s_28_port, PC_4out(27) => 
                           pc4_s_27_port, PC_4out(26) => pc4_s_26_port, 
                           PC_4out(25) => pc4_s_25_port, PC_4out(24) => 
                           pc4_s_24_port, PC_4out(23) => pc4_s_23_port, 
                           PC_4out(22) => pc4_s_22_port, PC_4out(21) => 
                           pc4_s_21_port, PC_4out(20) => pc4_s_20_port, 
                           PC_4out(19) => pc4_s_19_port, PC_4out(18) => 
                           pc4_s_18_port, PC_4out(17) => pc4_s_17_port, 
                           PC_4out(16) => pc4_s_16_port, PC_4out(15) => 
                           pc4_s_15_port, PC_4out(14) => pc4_s_14_port, 
                           PC_4out(13) => pc4_s_13_port, PC_4out(12) => 
                           pc4_s_12_port, PC_4out(11) => pc4_s_11_port, 
                           PC_4out(10) => pc4_s_10_port, PC_4out(9) => 
                           pc4_s_9_port, PC_4out(8) => pc4_s_8_port, PC_4out(7)
                           => pc4_s_7_port, PC_4out(6) => pc4_s_6_port, 
                           PC_4out(5) => pc4_s_5_port, PC_4out(4) => 
                           pc4_s_4_port, PC_4out(3) => pc4_s_3_port, PC_4out(2)
                           => pc4_s_2_port, PC_4out(1) => pc4_s_1_port, 
                           PC_4out(0) => pc4_s_0_port);
   D_STAGE : DU_N32 port map( J_EN => J_EN, WR_EN => RF_WE, A_EN => RegA_EN, 
                           B_EN => RegB_EN, IMM_EN => RegIMM_EN, RT_EN => 
                           RT_REG_EN, is_R_type => IS_R_TYPE, BR_EN => 
                           branch_taken_port, clk => CLK, rst => RST, 
                           NPC_IN(31) => npc_reg1_s_31_port, NPC_IN(30) => 
                           npc_reg1_s_30_port, NPC_IN(29) => npc_reg1_s_29_port
                           , NPC_IN(28) => npc_reg1_s_28_port, NPC_IN(27) => 
                           npc_reg1_s_27_port, NPC_IN(26) => npc_reg1_s_26_port
                           , NPC_IN(25) => npc_reg1_s_25_port, NPC_IN(24) => 
                           npc_reg1_s_24_port, NPC_IN(23) => npc_reg1_s_23_port
                           , NPC_IN(22) => npc_reg1_s_22_port, NPC_IN(21) => 
                           npc_reg1_s_21_port, NPC_IN(20) => npc_reg1_s_20_port
                           , NPC_IN(19) => npc_reg1_s_19_port, NPC_IN(18) => 
                           npc_reg1_s_18_port, NPC_IN(17) => npc_reg1_s_17_port
                           , NPC_IN(16) => npc_reg1_s_16_port, NPC_IN(15) => 
                           npc_reg1_s_15_port, NPC_IN(14) => npc_reg1_s_14_port
                           , NPC_IN(13) => npc_reg1_s_13_port, NPC_IN(12) => 
                           npc_reg1_s_12_port, NPC_IN(11) => npc_reg1_s_11_port
                           , NPC_IN(10) => npc_reg1_s_10_port, NPC_IN(9) => 
                           npc_reg1_s_9_port, NPC_IN(8) => npc_reg1_s_8_port, 
                           NPC_IN(7) => npc_reg1_s_7_port, NPC_IN(6) => 
                           npc_reg1_s_6_port, NPC_IN(5) => npc_reg1_s_5_port, 
                           NPC_IN(4) => npc_reg1_s_4_port, NPC_IN(3) => 
                           npc_reg1_s_3_port, NPC_IN(2) => npc_reg1_s_2_port, 
                           NPC_IN(1) => npc_reg1_s_1_port, NPC_IN(0) => 
                           npc_reg1_s_0_port, IR(31) => IR_31_port, IR(30) => 
                           IR_30_port, IR(29) => IR_29_port, IR(28) => 
                           IR_28_port, IR(27) => IR_27_port, IR(26) => 
                           IR_26_port, IR(25) => IR_25_port, IR(24) => 
                           IR_24_port, IR(23) => IR_23_port, IR(22) => 
                           IR_22_port, IR(21) => IR_21_port, IR(20) => 
                           IR_20_port, IR(19) => IR_19_port, IR(18) => 
                           IR_18_port, IR(17) => IR_17_port, IR(16) => 
                           IR_16_port, IR(15) => IR_15_port, IR(14) => 
                           IR_14_port, IR(13) => IR_13_port, IR(12) => 
                           IR_12_port, IR(11) => IR_11_port, IR(10) => 
                           IR_10_port, IR(9) => IR_9_port, IR(8) => IR_8_port, 
                           IR(7) => IR_7_port, IR(6) => IR_6_port, IR(5) => 
                           IR_5_port, IR(4) => IR_4_port, IR(3) => IR_3_port, 
                           IR(2) => IR_2_port, IR(1) => IR_1_port, IR(0) => 
                           IR_0_port, DATAIN(31) => wb_data_s_31_port, 
                           DATAIN(30) => wb_data_s_30_port, DATAIN(29) => 
                           wb_data_s_29_port, DATAIN(28) => wb_data_s_28_port, 
                           DATAIN(27) => wb_data_s_27_port, DATAIN(26) => 
                           wb_data_s_26_port, DATAIN(25) => wb_data_s_25_port, 
                           DATAIN(24) => wb_data_s_24_port, DATAIN(23) => 
                           wb_data_s_23_port, DATAIN(22) => wb_data_s_22_port, 
                           DATAIN(21) => wb_data_s_21_port, DATAIN(20) => 
                           wb_data_s_20_port, DATAIN(19) => wb_data_s_19_port, 
                           DATAIN(18) => wb_data_s_18_port, DATAIN(17) => 
                           wb_data_s_17_port, DATAIN(16) => wb_data_s_16_port, 
                           DATAIN(15) => wb_data_s_15_port, DATAIN(14) => 
                           wb_data_s_14_port, DATAIN(13) => wb_data_s_13_port, 
                           DATAIN(12) => wb_data_s_12_port, DATAIN(11) => 
                           wb_data_s_11_port, DATAIN(10) => wb_data_s_10_port, 
                           DATAIN(9) => wb_data_s_9_port, DATAIN(8) => 
                           wb_data_s_8_port, DATAIN(7) => wb_data_s_7_port, 
                           DATAIN(6) => wb_data_s_6_port, DATAIN(5) => 
                           wb_data_s_5_port, DATAIN(4) => wb_data_s_4_port, 
                           DATAIN(3) => wb_data_s_3_port, DATAIN(2) => 
                           wb_data_s_2_port, DATAIN(1) => wb_data_s_1_port, 
                           DATAIN(0) => wb_data_s_0_port, ADDR_IN(31) => 
                           wb_addr_s_31_port, ADDR_IN(30) => wb_addr_s_30_port,
                           ADDR_IN(29) => wb_addr_s_29_port, ADDR_IN(28) => 
                           wb_addr_s_28_port, ADDR_IN(27) => wb_addr_s_27_port,
                           ADDR_IN(26) => wb_addr_s_26_port, ADDR_IN(25) => 
                           wb_addr_s_25_port, ADDR_IN(24) => wb_addr_s_24_port,
                           ADDR_IN(23) => wb_addr_s_23_port, ADDR_IN(22) => 
                           wb_addr_s_22_port, ADDR_IN(21) => wb_addr_s_21_port,
                           ADDR_IN(20) => wb_addr_s_20_port, ADDR_IN(19) => 
                           wb_addr_s_19_port, ADDR_IN(18) => wb_addr_s_18_port,
                           ADDR_IN(17) => wb_addr_s_17_port, ADDR_IN(16) => 
                           wb_addr_s_16_port, ADDR_IN(15) => wb_addr_s_15_port,
                           ADDR_IN(14) => wb_addr_s_14_port, ADDR_IN(13) => 
                           wb_addr_s_13_port, ADDR_IN(12) => wb_addr_s_12_port,
                           ADDR_IN(11) => wb_addr_s_11_port, ADDR_IN(10) => 
                           wb_addr_s_10_port, ADDR_IN(9) => wb_addr_s_9_port, 
                           ADDR_IN(8) => wb_addr_s_8_port, ADDR_IN(7) => 
                           wb_addr_s_7_port, ADDR_IN(6) => wb_addr_s_6_port, 
                           ADDR_IN(5) => wb_addr_s_5_port, ADDR_IN(4) => 
                           wb_addr_s_4_port, ADDR_IN(3) => wb_addr_s_3_port, 
                           ADDR_IN(2) => wb_addr_s_2_port, ADDR_IN(1) => 
                           wb_addr_s_1_port, ADDR_IN(0) => wb_addr_s_0_port, 
                           BTA_OR_NPC(31) => b_addr_s_31_port, BTA_OR_NPC(30) 
                           => b_addr_s_30_port, BTA_OR_NPC(29) => 
                           b_addr_s_29_port, BTA_OR_NPC(28) => b_addr_s_28_port
                           , BTA_OR_NPC(27) => b_addr_s_27_port, BTA_OR_NPC(26)
                           => b_addr_s_26_port, BTA_OR_NPC(25) => 
                           b_addr_s_25_port, BTA_OR_NPC(24) => b_addr_s_24_port
                           , BTA_OR_NPC(23) => b_addr_s_23_port, BTA_OR_NPC(22)
                           => b_addr_s_22_port, BTA_OR_NPC(21) => 
                           b_addr_s_21_port, BTA_OR_NPC(20) => b_addr_s_20_port
                           , BTA_OR_NPC(19) => b_addr_s_19_port, BTA_OR_NPC(18)
                           => b_addr_s_18_port, BTA_OR_NPC(17) => 
                           b_addr_s_17_port, BTA_OR_NPC(16) => b_addr_s_16_port
                           , BTA_OR_NPC(15) => b_addr_s_15_port, BTA_OR_NPC(14)
                           => b_addr_s_14_port, BTA_OR_NPC(13) => 
                           b_addr_s_13_port, BTA_OR_NPC(12) => b_addr_s_12_port
                           , BTA_OR_NPC(11) => b_addr_s_11_port, BTA_OR_NPC(10)
                           => b_addr_s_10_port, BTA_OR_NPC(9) => 
                           b_addr_s_9_port, BTA_OR_NPC(8) => b_addr_s_8_port, 
                           BTA_OR_NPC(7) => b_addr_s_7_port, BTA_OR_NPC(6) => 
                           b_addr_s_6_port, BTA_OR_NPC(5) => b_addr_s_5_port, 
                           BTA_OR_NPC(4) => b_addr_s_4_port, BTA_OR_NPC(3) => 
                           b_addr_s_3_port, BTA_OR_NPC(2) => b_addr_s_2_port, 
                           BTA_OR_NPC(1) => b_addr_s_1_port, BTA_OR_NPC(0) => 
                           b_addr_s_0_port, A(31) => a_reg_s_31_port, A(30) => 
                           a_reg_s_30_port, A(29) => a_reg_s_29_port, A(28) => 
                           a_reg_s_28_port, A(27) => a_reg_s_27_port, A(26) => 
                           a_reg_s_26_port, A(25) => a_reg_s_25_port, A(24) => 
                           a_reg_s_24_port, A(23) => a_reg_s_23_port, A(22) => 
                           a_reg_s_22_port, A(21) => a_reg_s_21_port, A(20) => 
                           a_reg_s_20_port, A(19) => a_reg_s_19_port, A(18) => 
                           a_reg_s_18_port, A(17) => a_reg_s_17_port, A(16) => 
                           a_reg_s_16_port, A(15) => a_reg_s_15_port, A(14) => 
                           a_reg_s_14_port, A(13) => a_reg_s_13_port, A(12) => 
                           a_reg_s_12_port, A(11) => a_reg_s_11_port, A(10) => 
                           a_reg_s_10_port, A(9) => a_reg_s_9_port, A(8) => 
                           a_reg_s_8_port, A(7) => a_reg_s_7_port, A(6) => 
                           a_reg_s_6_port, A(5) => a_reg_s_5_port, A(4) => 
                           a_reg_s_4_port, A(3) => a_reg_s_3_port, A(2) => 
                           a_reg_s_2_port, A(1) => a_reg_s_1_port, A(0) => 
                           a_reg_s_0_port, B(31) => b_reg_s_31_port, B(30) => 
                           b_reg_s_30_port, B(29) => b_reg_s_29_port, B(28) => 
                           b_reg_s_28_port, B(27) => b_reg_s_27_port, B(26) => 
                           b_reg_s_26_port, B(25) => b_reg_s_25_port, B(24) => 
                           b_reg_s_24_port, B(23) => b_reg_s_23_port, B(22) => 
                           b_reg_s_22_port, B(21) => b_reg_s_21_port, B(20) => 
                           b_reg_s_20_port, B(19) => b_reg_s_19_port, B(18) => 
                           b_reg_s_18_port, B(17) => b_reg_s_17_port, B(16) => 
                           b_reg_s_16_port, B(15) => b_reg_s_15_port, B(14) => 
                           b_reg_s_14_port, B(13) => b_reg_s_13_port, B(12) => 
                           b_reg_s_12_port, B(11) => b_reg_s_11_port, B(10) => 
                           b_reg_s_10_port, B(9) => b_reg_s_9_port, B(8) => 
                           b_reg_s_8_port, B(7) => b_reg_s_7_port, B(6) => 
                           b_reg_s_6_port, B(5) => b_reg_s_5_port, B(4) => 
                           b_reg_s_4_port, B(3) => b_reg_s_3_port, B(2) => 
                           b_reg_s_2_port, B(1) => b_reg_s_1_port, B(0) => 
                           b_reg_s_0_port, IMM(31) => imm_reg_s_31_port, 
                           IMM(30) => imm_reg_s_30_port, IMM(29) => 
                           imm_reg_s_29_port, IMM(28) => imm_reg_s_28_port, 
                           IMM(27) => imm_reg_s_27_port, IMM(26) => 
                           imm_reg_s_26_port, IMM(25) => imm_reg_s_25_port, 
                           IMM(24) => imm_reg_s_24_port, IMM(23) => 
                           imm_reg_s_23_port, IMM(22) => imm_reg_s_22_port, 
                           IMM(21) => imm_reg_s_21_port, IMM(20) => 
                           imm_reg_s_20_port, IMM(19) => imm_reg_s_19_port, 
                           IMM(18) => imm_reg_s_18_port, IMM(17) => 
                           imm_reg_s_17_port, IMM(16) => imm_reg_s_16_port, 
                           IMM(15) => imm_reg_s_15_port, IMM(14) => 
                           imm_reg_s_14_port, IMM(13) => imm_reg_s_13_port, 
                           IMM(12) => imm_reg_s_12_port, IMM(11) => 
                           imm_reg_s_11_port, IMM(10) => imm_reg_s_10_port, 
                           IMM(9) => imm_reg_s_9_port, IMM(8) => 
                           imm_reg_s_8_port, IMM(7) => imm_reg_s_7_port, IMM(6)
                           => imm_reg_s_6_port, IMM(5) => imm_reg_s_5_port, 
                           IMM(4) => imm_reg_s_4_port, IMM(3) => 
                           imm_reg_s_3_port, IMM(2) => imm_reg_s_2_port, IMM(1)
                           => imm_reg_s_1_port, IMM(0) => imm_reg_s_0_port, 
                           RT_OUT(31) => rt_reg1_s_31_port, RT_OUT(30) => 
                           rt_reg1_s_30_port, RT_OUT(29) => rt_reg1_s_29_port, 
                           RT_OUT(28) => rt_reg1_s_28_port, RT_OUT(27) => 
                           rt_reg1_s_27_port, RT_OUT(26) => rt_reg1_s_26_port, 
                           RT_OUT(25) => rt_reg1_s_25_port, RT_OUT(24) => 
                           rt_reg1_s_24_port, RT_OUT(23) => rt_reg1_s_23_port, 
                           RT_OUT(22) => rt_reg1_s_22_port, RT_OUT(21) => 
                           rt_reg1_s_21_port, RT_OUT(20) => rt_reg1_s_20_port, 
                           RT_OUT(19) => rt_reg1_s_19_port, RT_OUT(18) => 
                           rt_reg1_s_18_port, RT_OUT(17) => rt_reg1_s_17_port, 
                           RT_OUT(16) => rt_reg1_s_16_port, RT_OUT(15) => 
                           rt_reg1_s_15_port, RT_OUT(14) => rt_reg1_s_14_port, 
                           RT_OUT(13) => rt_reg1_s_13_port, RT_OUT(12) => 
                           rt_reg1_s_12_port, RT_OUT(11) => rt_reg1_s_11_port, 
                           RT_OUT(10) => rt_reg1_s_10_port, RT_OUT(9) => 
                           rt_reg1_s_9_port, RT_OUT(8) => rt_reg1_s_8_port, 
                           RT_OUT(7) => rt_reg1_s_7_port, RT_OUT(6) => 
                           rt_reg1_s_6_port, RT_OUT(5) => rt_reg1_s_5_port, 
                           RT_OUT(4) => rt_reg1_s_4_port, RT_OUT(3) => 
                           rt_reg1_s_3_port, RT_OUT(2) => rt_reg1_s_2_port, 
                           RT_OUT(1) => rt_reg1_s_1_port, RT_OUT(0) => 
                           rt_reg1_s_0_port, NPC_OUT(31) => npc_reg2_s_31_port,
                           NPC_OUT(30) => npc_reg2_s_30_port, NPC_OUT(29) => 
                           npc_reg2_s_29_port, NPC_OUT(28) => 
                           npc_reg2_s_28_port, NPC_OUT(27) => 
                           npc_reg2_s_27_port, NPC_OUT(26) => 
                           npc_reg2_s_26_port, NPC_OUT(25) => 
                           npc_reg2_s_25_port, NPC_OUT(24) => 
                           npc_reg2_s_24_port, NPC_OUT(23) => 
                           npc_reg2_s_23_port, NPC_OUT(22) => 
                           npc_reg2_s_22_port, NPC_OUT(21) => 
                           npc_reg2_s_21_port, NPC_OUT(20) => 
                           npc_reg2_s_20_port, NPC_OUT(19) => 
                           npc_reg2_s_19_port, NPC_OUT(18) => 
                           npc_reg2_s_18_port, NPC_OUT(17) => 
                           npc_reg2_s_17_port, NPC_OUT(16) => 
                           npc_reg2_s_16_port, NPC_OUT(15) => 
                           npc_reg2_s_15_port, NPC_OUT(14) => 
                           npc_reg2_s_14_port, NPC_OUT(13) => 
                           npc_reg2_s_13_port, NPC_OUT(12) => 
                           npc_reg2_s_12_port, NPC_OUT(11) => 
                           npc_reg2_s_11_port, NPC_OUT(10) => 
                           npc_reg2_s_10_port, NPC_OUT(9) => npc_reg2_s_9_port,
                           NPC_OUT(8) => npc_reg2_s_8_port, NPC_OUT(7) => 
                           npc_reg2_s_7_port, NPC_OUT(6) => npc_reg2_s_6_port, 
                           NPC_OUT(5) => npc_reg2_s_5_port, NPC_OUT(4) => 
                           npc_reg2_s_4_port, NPC_OUT(3) => npc_reg2_s_3_port, 
                           NPC_OUT(2) => npc_reg2_s_2_port, NPC_OUT(1) => 
                           npc_reg2_s_1_port, NPC_OUT(0) => npc_reg2_s_0_port, 
                           PC_NXT(31) => pc_nxt_s_31_port, PC_NXT(30) => 
                           pc_nxt_s_30_port, PC_NXT(29) => pc_nxt_s_29_port, 
                           PC_NXT(28) => pc_nxt_s_28_port, PC_NXT(27) => 
                           pc_nxt_s_27_port, PC_NXT(26) => pc_nxt_s_26_port, 
                           PC_NXT(25) => pc_nxt_s_25_port, PC_NXT(24) => 
                           pc_nxt_s_24_port, PC_NXT(23) => pc_nxt_s_23_port, 
                           PC_NXT(22) => pc_nxt_s_22_port, PC_NXT(21) => 
                           pc_nxt_s_21_port, PC_NXT(20) => pc_nxt_s_20_port, 
                           PC_NXT(19) => pc_nxt_s_19_port, PC_NXT(18) => 
                           pc_nxt_s_18_port, PC_NXT(17) => pc_nxt_s_17_port, 
                           PC_NXT(16) => pc_nxt_s_16_port, PC_NXT(15) => 
                           pc_nxt_s_15_port, PC_NXT(14) => pc_nxt_s_14_port, 
                           PC_NXT(13) => pc_nxt_s_13_port, PC_NXT(12) => 
                           pc_nxt_s_12_port, PC_NXT(11) => pc_nxt_s_11_port, 
                           PC_NXT(10) => pc_nxt_s_10_port, PC_NXT(9) => 
                           pc_nxt_s_9_port, PC_NXT(8) => pc_nxt_s_8_port, 
                           PC_NXT(7) => pc_nxt_s_7_port, PC_NXT(6) => 
                           pc_nxt_s_6_port, PC_NXT(5) => pc_nxt_s_5_port, 
                           PC_NXT(4) => pc_nxt_s_4_port, PC_NXT(3) => 
                           pc_nxt_s_3_port, PC_NXT(2) => pc_nxt_s_2_port, 
                           PC_NXT(1) => pc_nxt_s_1_port, PC_NXT(0) => 
                           pc_nxt_s_0_port);
   EX_STAGE : EXU_N32 port map( CLK => CLK, RST => RST, MUXA_SEL => MUXA_SEL, 
                           MUXB_SEL => MUXB_SEL, ZERO_EN => BRANCH_EN, ZERO_SEL
                           => BEQZ_OR_BNEZ, ALUOUT_EN => ALU_OUTREG_EN, 
                           SHIFT2_EN => SH2_EN, ALU_FUNC(0) => ALU_FUNC(0), 
                           ALU_FUNC(1) => ALU_FUNC(1), ALU_FUNC(2) => 
                           ALU_FUNC(2), ALU_FUNC(3) => ALU_FUNC(3), NPC_REG(31)
                           => npc_reg2_s_31_port, NPC_REG(30) => 
                           npc_reg2_s_30_port, NPC_REG(29) => 
                           npc_reg2_s_29_port, NPC_REG(28) => 
                           npc_reg2_s_28_port, NPC_REG(27) => 
                           npc_reg2_s_27_port, NPC_REG(26) => 
                           npc_reg2_s_26_port, NPC_REG(25) => 
                           npc_reg2_s_25_port, NPC_REG(24) => 
                           npc_reg2_s_24_port, NPC_REG(23) => 
                           npc_reg2_s_23_port, NPC_REG(22) => 
                           npc_reg2_s_22_port, NPC_REG(21) => 
                           npc_reg2_s_21_port, NPC_REG(20) => 
                           npc_reg2_s_20_port, NPC_REG(19) => 
                           npc_reg2_s_19_port, NPC_REG(18) => 
                           npc_reg2_s_18_port, NPC_REG(17) => 
                           npc_reg2_s_17_port, NPC_REG(16) => 
                           npc_reg2_s_16_port, NPC_REG(15) => 
                           npc_reg2_s_15_port, NPC_REG(14) => 
                           npc_reg2_s_14_port, NPC_REG(13) => 
                           npc_reg2_s_13_port, NPC_REG(12) => 
                           npc_reg2_s_12_port, NPC_REG(11) => 
                           npc_reg2_s_11_port, NPC_REG(10) => 
                           npc_reg2_s_10_port, NPC_REG(9) => npc_reg2_s_9_port,
                           NPC_REG(8) => npc_reg2_s_8_port, NPC_REG(7) => 
                           npc_reg2_s_7_port, NPC_REG(6) => npc_reg2_s_6_port, 
                           NPC_REG(5) => npc_reg2_s_5_port, NPC_REG(4) => 
                           npc_reg2_s_4_port, NPC_REG(3) => npc_reg2_s_3_port, 
                           NPC_REG(2) => npc_reg2_s_2_port, NPC_REG(1) => 
                           npc_reg2_s_1_port, NPC_REG(0) => npc_reg2_s_0_port, 
                           A_REG(31) => a_reg_s_31_port, A_REG(30) => 
                           a_reg_s_30_port, A_REG(29) => a_reg_s_29_port, 
                           A_REG(28) => a_reg_s_28_port, A_REG(27) => 
                           a_reg_s_27_port, A_REG(26) => a_reg_s_26_port, 
                           A_REG(25) => a_reg_s_25_port, A_REG(24) => 
                           a_reg_s_24_port, A_REG(23) => a_reg_s_23_port, 
                           A_REG(22) => a_reg_s_22_port, A_REG(21) => 
                           a_reg_s_21_port, A_REG(20) => a_reg_s_20_port, 
                           A_REG(19) => a_reg_s_19_port, A_REG(18) => 
                           a_reg_s_18_port, A_REG(17) => a_reg_s_17_port, 
                           A_REG(16) => a_reg_s_16_port, A_REG(15) => 
                           a_reg_s_15_port, A_REG(14) => a_reg_s_14_port, 
                           A_REG(13) => a_reg_s_13_port, A_REG(12) => 
                           a_reg_s_12_port, A_REG(11) => a_reg_s_11_port, 
                           A_REG(10) => a_reg_s_10_port, A_REG(9) => 
                           a_reg_s_9_port, A_REG(8) => a_reg_s_8_port, A_REG(7)
                           => a_reg_s_7_port, A_REG(6) => a_reg_s_6_port, 
                           A_REG(5) => a_reg_s_5_port, A_REG(4) => 
                           a_reg_s_4_port, A_REG(3) => a_reg_s_3_port, A_REG(2)
                           => a_reg_s_2_port, A_REG(1) => a_reg_s_1_port, 
                           A_REG(0) => a_reg_s_0_port, B_REG(31) => 
                           b_reg_s_31_port, B_REG(30) => b_reg_s_30_port, 
                           B_REG(29) => b_reg_s_29_port, B_REG(28) => 
                           b_reg_s_28_port, B_REG(27) => b_reg_s_27_port, 
                           B_REG(26) => b_reg_s_26_port, B_REG(25) => 
                           b_reg_s_25_port, B_REG(24) => b_reg_s_24_port, 
                           B_REG(23) => b_reg_s_23_port, B_REG(22) => 
                           b_reg_s_22_port, B_REG(21) => b_reg_s_21_port, 
                           B_REG(20) => b_reg_s_20_port, B_REG(19) => 
                           b_reg_s_19_port, B_REG(18) => b_reg_s_18_port, 
                           B_REG(17) => b_reg_s_17_port, B_REG(16) => 
                           b_reg_s_16_port, B_REG(15) => b_reg_s_15_port, 
                           B_REG(14) => b_reg_s_14_port, B_REG(13) => 
                           b_reg_s_13_port, B_REG(12) => b_reg_s_12_port, 
                           B_REG(11) => b_reg_s_11_port, B_REG(10) => 
                           b_reg_s_10_port, B_REG(9) => b_reg_s_9_port, 
                           B_REG(8) => b_reg_s_8_port, B_REG(7) => 
                           b_reg_s_7_port, B_REG(6) => b_reg_s_6_port, B_REG(5)
                           => b_reg_s_5_port, B_REG(4) => b_reg_s_4_port, 
                           B_REG(3) => b_reg_s_3_port, B_REG(2) => 
                           b_reg_s_2_port, B_REG(1) => b_reg_s_1_port, B_REG(0)
                           => b_reg_s_0_port, RT_REG(31) => rt_reg1_s_31_port, 
                           RT_REG(30) => rt_reg1_s_30_port, RT_REG(29) => 
                           rt_reg1_s_29_port, RT_REG(28) => rt_reg1_s_28_port, 
                           RT_REG(27) => rt_reg1_s_27_port, RT_REG(26) => 
                           rt_reg1_s_26_port, RT_REG(25) => rt_reg1_s_25_port, 
                           RT_REG(24) => rt_reg1_s_24_port, RT_REG(23) => 
                           rt_reg1_s_23_port, RT_REG(22) => rt_reg1_s_22_port, 
                           RT_REG(21) => rt_reg1_s_21_port, RT_REG(20) => 
                           rt_reg1_s_20_port, RT_REG(19) => rt_reg1_s_19_port, 
                           RT_REG(18) => rt_reg1_s_18_port, RT_REG(17) => 
                           rt_reg1_s_17_port, RT_REG(16) => rt_reg1_s_16_port, 
                           RT_REG(15) => rt_reg1_s_15_port, RT_REG(14) => 
                           rt_reg1_s_14_port, RT_REG(13) => rt_reg1_s_13_port, 
                           RT_REG(12) => rt_reg1_s_12_port, RT_REG(11) => 
                           rt_reg1_s_11_port, RT_REG(10) => rt_reg1_s_10_port, 
                           RT_REG(9) => rt_reg1_s_9_port, RT_REG(8) => 
                           rt_reg1_s_8_port, RT_REG(7) => rt_reg1_s_7_port, 
                           RT_REG(6) => rt_reg1_s_6_port, RT_REG(5) => 
                           rt_reg1_s_5_port, RT_REG(4) => rt_reg1_s_4_port, 
                           RT_REG(3) => rt_reg1_s_3_port, RT_REG(2) => 
                           rt_reg1_s_2_port, RT_REG(1) => rt_reg1_s_1_port, 
                           RT_REG(0) => rt_reg1_s_0_port, IMM_REG(31) => 
                           imm_reg_s_31_port, IMM_REG(30) => imm_reg_s_30_port,
                           IMM_REG(29) => imm_reg_s_29_port, IMM_REG(28) => 
                           imm_reg_s_28_port, IMM_REG(27) => imm_reg_s_27_port,
                           IMM_REG(26) => imm_reg_s_26_port, IMM_REG(25) => 
                           imm_reg_s_25_port, IMM_REG(24) => imm_reg_s_24_port,
                           IMM_REG(23) => imm_reg_s_23_port, IMM_REG(22) => 
                           imm_reg_s_22_port, IMM_REG(21) => imm_reg_s_21_port,
                           IMM_REG(20) => imm_reg_s_20_port, IMM_REG(19) => 
                           imm_reg_s_19_port, IMM_REG(18) => imm_reg_s_18_port,
                           IMM_REG(17) => imm_reg_s_17_port, IMM_REG(16) => 
                           imm_reg_s_16_port, IMM_REG(15) => imm_reg_s_15_port,
                           IMM_REG(14) => imm_reg_s_14_port, IMM_REG(13) => 
                           imm_reg_s_13_port, IMM_REG(12) => imm_reg_s_12_port,
                           IMM_REG(11) => imm_reg_s_11_port, IMM_REG(10) => 
                           imm_reg_s_10_port, IMM_REG(9) => imm_reg_s_9_port, 
                           IMM_REG(8) => imm_reg_s_8_port, IMM_REG(7) => 
                           imm_reg_s_7_port, IMM_REG(6) => imm_reg_s_6_port, 
                           IMM_REG(5) => imm_reg_s_5_port, IMM_REG(4) => 
                           imm_reg_s_4_port, IMM_REG(3) => imm_reg_s_3_port, 
                           IMM_REG(2) => imm_reg_s_2_port, IMM_REG(1) => 
                           imm_reg_s_1_port, IMM_REG(0) => imm_reg_s_0_port, 
                           PC_4(31) => pc4_s_31_port, PC_4(30) => pc4_s_30_port
                           , PC_4(29) => pc4_s_29_port, PC_4(28) => 
                           pc4_s_28_port, PC_4(27) => pc4_s_27_port, PC_4(26) 
                           => pc4_s_26_port, PC_4(25) => pc4_s_25_port, 
                           PC_4(24) => pc4_s_24_port, PC_4(23) => pc4_s_23_port
                           , PC_4(22) => pc4_s_22_port, PC_4(21) => 
                           pc4_s_21_port, PC_4(20) => pc4_s_20_port, PC_4(19) 
                           => pc4_s_19_port, PC_4(18) => pc4_s_18_port, 
                           PC_4(17) => pc4_s_17_port, PC_4(16) => pc4_s_16_port
                           , PC_4(15) => pc4_s_15_port, PC_4(14) => 
                           pc4_s_14_port, PC_4(13) => pc4_s_13_port, PC_4(12) 
                           => pc4_s_12_port, PC_4(11) => pc4_s_11_port, 
                           PC_4(10) => pc4_s_10_port, PC_4(9) => pc4_s_9_port, 
                           PC_4(8) => pc4_s_8_port, PC_4(7) => pc4_s_7_port, 
                           PC_4(6) => pc4_s_6_port, PC_4(5) => pc4_s_5_port, 
                           PC_4(4) => pc4_s_4_port, PC_4(3) => pc4_s_3_port, 
                           PC_4(2) => pc4_s_2_port, PC_4(1) => pc4_s_1_port, 
                           PC_4(0) => pc4_s_0_port, ZERO => branch_taken_port, 
                           BRANC_ADDR(31) => b_addr_s_31_port, BRANC_ADDR(30) 
                           => b_addr_s_30_port, BRANC_ADDR(29) => 
                           b_addr_s_29_port, BRANC_ADDR(28) => b_addr_s_28_port
                           , BRANC_ADDR(27) => b_addr_s_27_port, BRANC_ADDR(26)
                           => b_addr_s_26_port, BRANC_ADDR(25) => 
                           b_addr_s_25_port, BRANC_ADDR(24) => b_addr_s_24_port
                           , BRANC_ADDR(23) => b_addr_s_23_port, BRANC_ADDR(22)
                           => b_addr_s_22_port, BRANC_ADDR(21) => 
                           b_addr_s_21_port, BRANC_ADDR(20) => b_addr_s_20_port
                           , BRANC_ADDR(19) => b_addr_s_19_port, BRANC_ADDR(18)
                           => b_addr_s_18_port, BRANC_ADDR(17) => 
                           b_addr_s_17_port, BRANC_ADDR(16) => b_addr_s_16_port
                           , BRANC_ADDR(15) => b_addr_s_15_port, BRANC_ADDR(14)
                           => b_addr_s_14_port, BRANC_ADDR(13) => 
                           b_addr_s_13_port, BRANC_ADDR(12) => b_addr_s_12_port
                           , BRANC_ADDR(11) => b_addr_s_11_port, BRANC_ADDR(10)
                           => b_addr_s_10_port, BRANC_ADDR(9) => 
                           b_addr_s_9_port, BRANC_ADDR(8) => b_addr_s_8_port, 
                           BRANC_ADDR(7) => b_addr_s_7_port, BRANC_ADDR(6) => 
                           b_addr_s_6_port, BRANC_ADDR(5) => b_addr_s_5_port, 
                           BRANC_ADDR(4) => b_addr_s_4_port, BRANC_ADDR(3) => 
                           b_addr_s_3_port, BRANC_ADDR(2) => b_addr_s_2_port, 
                           BRANC_ADDR(1) => b_addr_s_1_port, BRANC_ADDR(0) => 
                           b_addr_s_0_port, ALU_OUT(31) => addr_to_DRAM_31_port
                           , ALU_OUT(30) => addr_to_DRAM_30_port, ALU_OUT(29) 
                           => addr_to_DRAM_29_port, ALU_OUT(28) => 
                           addr_to_DRAM_28_port, ALU_OUT(27) => 
                           addr_to_DRAM_27_port, ALU_OUT(26) => 
                           addr_to_DRAM_26_port, ALU_OUT(25) => 
                           addr_to_DRAM_25_port, ALU_OUT(24) => 
                           addr_to_DRAM_24_port, ALU_OUT(23) => 
                           addr_to_DRAM_23_port, ALU_OUT(22) => 
                           addr_to_DRAM_22_port, ALU_OUT(21) => 
                           addr_to_DRAM_21_port, ALU_OUT(20) => 
                           addr_to_DRAM_20_port, ALU_OUT(19) => 
                           addr_to_DRAM_19_port, ALU_OUT(18) => 
                           addr_to_DRAM_18_port, ALU_OUT(17) => 
                           addr_to_DRAM_17_port, ALU_OUT(16) => 
                           addr_to_DRAM_16_port, ALU_OUT(15) => 
                           addr_to_DRAM_15_port, ALU_OUT(14) => 
                           addr_to_DRAM_14_port, ALU_OUT(13) => 
                           addr_to_DRAM_13_port, ALU_OUT(12) => 
                           addr_to_DRAM_12_port, ALU_OUT(11) => 
                           addr_to_DRAM_11_port, ALU_OUT(10) => 
                           addr_to_DRAM_10_port, ALU_OUT(9) => 
                           addr_to_DRAM_9_port, ALU_OUT(8) => 
                           addr_to_DRAM_8_port, ALU_OUT(7) => 
                           addr_to_DRAM_7_port, ALU_OUT(6) => 
                           addr_to_DRAM_6_port, ALU_OUT(5) => 
                           addr_to_DRAM_5_port, ALU_OUT(4) => 
                           addr_to_DRAM_4_port, ALU_OUT(3) => 
                           addr_to_DRAM_3_port, ALU_OUT(2) => 
                           addr_to_DRAM_2_port, ALU_OUT(1) => 
                           addr_to_DRAM_1_port, ALU_OUT(0) => 
                           addr_to_DRAM_0_port, RT_REG_OUT(31) => 
                           data_to_DRAM_31_port, RT_REG_OUT(30) => 
                           data_to_DRAM_30_port, RT_REG_OUT(29) => 
                           data_to_DRAM_29_port, RT_REG_OUT(28) => 
                           data_to_DRAM_28_port, RT_REG_OUT(27) => 
                           data_to_DRAM_27_port, RT_REG_OUT(26) => 
                           data_to_DRAM_26_port, RT_REG_OUT(25) => 
                           data_to_DRAM_25_port, RT_REG_OUT(24) => 
                           data_to_DRAM_24_port, RT_REG_OUT(23) => 
                           data_to_DRAM_23_port, RT_REG_OUT(22) => 
                           data_to_DRAM_22_port, RT_REG_OUT(21) => 
                           data_to_DRAM_21_port, RT_REG_OUT(20) => 
                           data_to_DRAM_20_port, RT_REG_OUT(19) => 
                           data_to_DRAM_19_port, RT_REG_OUT(18) => 
                           data_to_DRAM_18_port, RT_REG_OUT(17) => 
                           data_to_DRAM_17_port, RT_REG_OUT(16) => 
                           data_to_DRAM_16_port, RT_REG_OUT(15) => 
                           data_to_DRAM_15_port, RT_REG_OUT(14) => 
                           data_to_DRAM_14_port, RT_REG_OUT(13) => 
                           data_to_DRAM_13_port, RT_REG_OUT(12) => 
                           data_to_DRAM_12_port, RT_REG_OUT(11) => 
                           data_to_DRAM_11_port, RT_REG_OUT(10) => 
                           data_to_DRAM_10_port, RT_REG_OUT(9) => 
                           data_to_DRAM_9_port, RT_REG_OUT(8) => 
                           data_to_DRAM_8_port, RT_REG_OUT(7) => 
                           data_to_DRAM_7_port, RT_REG_OUT(6) => 
                           data_to_DRAM_6_port, RT_REG_OUT(5) => 
                           data_to_DRAM_5_port, RT_REG_OUT(4) => 
                           data_to_DRAM_4_port, RT_REG_OUT(3) => 
                           data_to_DRAM_3_port, RT_REG_OUT(2) => 
                           data_to_DRAM_2_port, RT_REG_OUT(1) => 
                           data_to_DRAM_1_port, RT_REG_OUT(0) => 
                           data_to_DRAM_0_port, NPC_OUT(31) => 
                           npc_reg3_s_31_port, NPC_OUT(30) => 
                           npc_reg3_s_30_port, NPC_OUT(29) => 
                           npc_reg3_s_29_port, NPC_OUT(28) => 
                           npc_reg3_s_28_port, NPC_OUT(27) => 
                           npc_reg3_s_27_port, NPC_OUT(26) => 
                           npc_reg3_s_26_port, NPC_OUT(25) => 
                           npc_reg3_s_25_port, NPC_OUT(24) => 
                           npc_reg3_s_24_port, NPC_OUT(23) => 
                           npc_reg3_s_23_port, NPC_OUT(22) => 
                           npc_reg3_s_22_port, NPC_OUT(21) => 
                           npc_reg3_s_21_port, NPC_OUT(20) => 
                           npc_reg3_s_20_port, NPC_OUT(19) => 
                           npc_reg3_s_19_port, NPC_OUT(18) => 
                           npc_reg3_s_18_port, NPC_OUT(17) => 
                           npc_reg3_s_17_port, NPC_OUT(16) => 
                           npc_reg3_s_16_port, NPC_OUT(15) => 
                           npc_reg3_s_15_port, NPC_OUT(14) => 
                           npc_reg3_s_14_port, NPC_OUT(13) => 
                           npc_reg3_s_13_port, NPC_OUT(12) => 
                           npc_reg3_s_12_port, NPC_OUT(11) => 
                           npc_reg3_s_11_port, NPC_OUT(10) => 
                           npc_reg3_s_10_port, NPC_OUT(9) => npc_reg3_s_9_port,
                           NPC_OUT(8) => npc_reg3_s_8_port, NPC_OUT(7) => 
                           npc_reg3_s_7_port, NPC_OUT(6) => npc_reg3_s_6_port, 
                           NPC_OUT(5) => npc_reg3_s_5_port, NPC_OUT(4) => 
                           npc_reg3_s_4_port, NPC_OUT(3) => npc_reg3_s_3_port, 
                           NPC_OUT(2) => npc_reg3_s_2_port, NPC_OUT(1) => 
                           npc_reg3_s_1_port, NPC_OUT(0) => npc_reg3_s_0_port);
   MEM_STAGE : MU_N32 port map( CLK => CLK, RST => RST, LMD_EN => LMD_EN, 
                           ALU_RESULT(31) => addr_to_DRAM_31_port, 
                           ALU_RESULT(30) => addr_to_DRAM_30_port, 
                           ALU_RESULT(29) => addr_to_DRAM_29_port, 
                           ALU_RESULT(28) => addr_to_DRAM_28_port, 
                           ALU_RESULT(27) => addr_to_DRAM_27_port, 
                           ALU_RESULT(26) => addr_to_DRAM_26_port, 
                           ALU_RESULT(25) => addr_to_DRAM_25_port, 
                           ALU_RESULT(24) => addr_to_DRAM_24_port, 
                           ALU_RESULT(23) => addr_to_DRAM_23_port, 
                           ALU_RESULT(22) => addr_to_DRAM_22_port, 
                           ALU_RESULT(21) => addr_to_DRAM_21_port, 
                           ALU_RESULT(20) => addr_to_DRAM_20_port, 
                           ALU_RESULT(19) => addr_to_DRAM_19_port, 
                           ALU_RESULT(18) => addr_to_DRAM_18_port, 
                           ALU_RESULT(17) => addr_to_DRAM_17_port, 
                           ALU_RESULT(16) => addr_to_DRAM_16_port, 
                           ALU_RESULT(15) => addr_to_DRAM_15_port, 
                           ALU_RESULT(14) => addr_to_DRAM_14_port, 
                           ALU_RESULT(13) => addr_to_DRAM_13_port, 
                           ALU_RESULT(12) => addr_to_DRAM_12_port, 
                           ALU_RESULT(11) => addr_to_DRAM_11_port, 
                           ALU_RESULT(10) => addr_to_DRAM_10_port, 
                           ALU_RESULT(9) => addr_to_DRAM_9_port, ALU_RESULT(8) 
                           => addr_to_DRAM_8_port, ALU_RESULT(7) => 
                           addr_to_DRAM_7_port, ALU_RESULT(6) => 
                           addr_to_DRAM_6_port, ALU_RESULT(5) => 
                           addr_to_DRAM_5_port, ALU_RESULT(4) => 
                           addr_to_DRAM_4_port, ALU_RESULT(3) => 
                           addr_to_DRAM_3_port, ALU_RESULT(2) => 
                           addr_to_DRAM_2_port, ALU_RESULT(1) => 
                           addr_to_DRAM_1_port, ALU_RESULT(0) => 
                           addr_to_DRAM_0_port, RT_REG_in(31) => 
                           data_to_DRAM_31_port, RT_REG_in(30) => 
                           data_to_DRAM_30_port, RT_REG_in(29) => 
                           data_to_DRAM_29_port, RT_REG_in(28) => 
                           data_to_DRAM_28_port, RT_REG_in(27) => 
                           data_to_DRAM_27_port, RT_REG_in(26) => 
                           data_to_DRAM_26_port, RT_REG_in(25) => 
                           data_to_DRAM_25_port, RT_REG_in(24) => 
                           data_to_DRAM_24_port, RT_REG_in(23) => 
                           data_to_DRAM_23_port, RT_REG_in(22) => 
                           data_to_DRAM_22_port, RT_REG_in(21) => 
                           data_to_DRAM_21_port, RT_REG_in(20) => 
                           data_to_DRAM_20_port, RT_REG_in(19) => 
                           data_to_DRAM_19_port, RT_REG_in(18) => 
                           data_to_DRAM_18_port, RT_REG_in(17) => 
                           data_to_DRAM_17_port, RT_REG_in(16) => 
                           data_to_DRAM_16_port, RT_REG_in(15) => 
                           data_to_DRAM_15_port, RT_REG_in(14) => 
                           data_to_DRAM_14_port, RT_REG_in(13) => 
                           data_to_DRAM_13_port, RT_REG_in(12) => 
                           data_to_DRAM_12_port, RT_REG_in(11) => 
                           data_to_DRAM_11_port, RT_REG_in(10) => 
                           data_to_DRAM_10_port, RT_REG_in(9) => 
                           data_to_DRAM_9_port, RT_REG_in(8) => 
                           data_to_DRAM_8_port, RT_REG_in(7) => 
                           data_to_DRAM_7_port, RT_REG_in(6) => 
                           data_to_DRAM_6_port, RT_REG_in(5) => 
                           data_to_DRAM_5_port, RT_REG_in(4) => 
                           data_to_DRAM_4_port, RT_REG_in(3) => 
                           data_to_DRAM_3_port, RT_REG_in(2) => 
                           data_to_DRAM_2_port, RT_REG_in(1) => 
                           data_to_DRAM_1_port, RT_REG_in(0) => 
                           data_to_DRAM_0_port, NPC_REG_in(31) => 
                           npc_reg3_s_31_port, NPC_REG_in(30) => 
                           npc_reg3_s_30_port, NPC_REG_in(29) => 
                           npc_reg3_s_29_port, NPC_REG_in(28) => 
                           npc_reg3_s_28_port, NPC_REG_in(27) => 
                           npc_reg3_s_27_port, NPC_REG_in(26) => 
                           npc_reg3_s_26_port, NPC_REG_in(25) => 
                           npc_reg3_s_25_port, NPC_REG_in(24) => 
                           npc_reg3_s_24_port, NPC_REG_in(23) => 
                           npc_reg3_s_23_port, NPC_REG_in(22) => 
                           npc_reg3_s_22_port, NPC_REG_in(21) => 
                           npc_reg3_s_21_port, NPC_REG_in(20) => 
                           npc_reg3_s_20_port, NPC_REG_in(19) => 
                           npc_reg3_s_19_port, NPC_REG_in(18) => 
                           npc_reg3_s_18_port, NPC_REG_in(17) => 
                           npc_reg3_s_17_port, NPC_REG_in(16) => 
                           npc_reg3_s_16_port, NPC_REG_in(15) => 
                           npc_reg3_s_15_port, NPC_REG_in(14) => 
                           npc_reg3_s_14_port, NPC_REG_in(13) => 
                           npc_reg3_s_13_port, NPC_REG_in(12) => 
                           npc_reg3_s_12_port, NPC_REG_in(11) => 
                           npc_reg3_s_11_port, NPC_REG_in(10) => 
                           npc_reg3_s_10_port, NPC_REG_in(9) => 
                           npc_reg3_s_9_port, NPC_REG_in(8) => 
                           npc_reg3_s_8_port, NPC_REG_in(7) => 
                           npc_reg3_s_7_port, NPC_REG_in(6) => 
                           npc_reg3_s_6_port, NPC_REG_in(5) => 
                           npc_reg3_s_5_port, NPC_REG_in(4) => 
                           npc_reg3_s_4_port, NPC_REG_in(3) => 
                           npc_reg3_s_3_port, NPC_REG_in(2) => 
                           npc_reg3_s_2_port, NPC_REG_in(1) => 
                           npc_reg3_s_1_port, NPC_REG_in(0) => 
                           npc_reg3_s_0_port, LMD_LATCH_in(31) => from_DRAM(31)
                           , LMD_LATCH_in(30) => from_DRAM(30), 
                           LMD_LATCH_in(29) => from_DRAM(29), LMD_LATCH_in(28) 
                           => from_DRAM(28), LMD_LATCH_in(27) => from_DRAM(27),
                           LMD_LATCH_in(26) => from_DRAM(26), LMD_LATCH_in(25) 
                           => from_DRAM(25), LMD_LATCH_in(24) => from_DRAM(24),
                           LMD_LATCH_in(23) => from_DRAM(23), LMD_LATCH_in(22) 
                           => from_DRAM(22), LMD_LATCH_in(21) => from_DRAM(21),
                           LMD_LATCH_in(20) => from_DRAM(20), LMD_LATCH_in(19) 
                           => from_DRAM(19), LMD_LATCH_in(18) => from_DRAM(18),
                           LMD_LATCH_in(17) => from_DRAM(17), LMD_LATCH_in(16) 
                           => from_DRAM(16), LMD_LATCH_in(15) => from_DRAM(15),
                           LMD_LATCH_in(14) => from_DRAM(14), LMD_LATCH_in(13) 
                           => from_DRAM(13), LMD_LATCH_in(12) => from_DRAM(12),
                           LMD_LATCH_in(11) => from_DRAM(11), LMD_LATCH_in(10) 
                           => from_DRAM(10), LMD_LATCH_in(9) => from_DRAM(9), 
                           LMD_LATCH_in(8) => from_DRAM(8), LMD_LATCH_in(7) => 
                           from_DRAM(7), LMD_LATCH_in(6) => from_DRAM(6), 
                           LMD_LATCH_in(5) => from_DRAM(5), LMD_LATCH_in(4) => 
                           from_DRAM(4), LMD_LATCH_in(3) => from_DRAM(3), 
                           LMD_LATCH_in(2) => from_DRAM(2), LMD_LATCH_in(1) => 
                           from_DRAM(1), LMD_LATCH_in(0) => from_DRAM(0), 
                           LMD_LATCH_out(31) => lmd_out_s_31_port, 
                           LMD_LATCH_out(30) => lmd_out_s_30_port, 
                           LMD_LATCH_out(29) => lmd_out_s_29_port, 
                           LMD_LATCH_out(28) => lmd_out_s_28_port, 
                           LMD_LATCH_out(27) => lmd_out_s_27_port, 
                           LMD_LATCH_out(26) => lmd_out_s_26_port, 
                           LMD_LATCH_out(25) => lmd_out_s_25_port, 
                           LMD_LATCH_out(24) => lmd_out_s_24_port, 
                           LMD_LATCH_out(23) => lmd_out_s_23_port, 
                           LMD_LATCH_out(22) => lmd_out_s_22_port, 
                           LMD_LATCH_out(21) => lmd_out_s_21_port, 
                           LMD_LATCH_out(20) => lmd_out_s_20_port, 
                           LMD_LATCH_out(19) => lmd_out_s_19_port, 
                           LMD_LATCH_out(18) => lmd_out_s_18_port, 
                           LMD_LATCH_out(17) => lmd_out_s_17_port, 
                           LMD_LATCH_out(16) => lmd_out_s_16_port, 
                           LMD_LATCH_out(15) => lmd_out_s_15_port, 
                           LMD_LATCH_out(14) => lmd_out_s_14_port, 
                           LMD_LATCH_out(13) => lmd_out_s_13_port, 
                           LMD_LATCH_out(12) => lmd_out_s_12_port, 
                           LMD_LATCH_out(11) => lmd_out_s_11_port, 
                           LMD_LATCH_out(10) => lmd_out_s_10_port, 
                           LMD_LATCH_out(9) => lmd_out_s_9_port, 
                           LMD_LATCH_out(8) => lmd_out_s_8_port, 
                           LMD_LATCH_out(7) => lmd_out_s_7_port, 
                           LMD_LATCH_out(6) => lmd_out_s_6_port, 
                           LMD_LATCH_out(5) => lmd_out_s_5_port, 
                           LMD_LATCH_out(4) => lmd_out_s_4_port, 
                           LMD_LATCH_out(3) => lmd_out_s_3_port, 
                           LMD_LATCH_out(2) => lmd_out_s_2_port, 
                           LMD_LATCH_out(1) => lmd_out_s_1_port, 
                           LMD_LATCH_out(0) => lmd_out_s_0_port, 
                           ALU_REG_out(31) => alu_out2_s_31_port, 
                           ALU_REG_out(30) => alu_out2_s_30_port, 
                           ALU_REG_out(29) => alu_out2_s_29_port, 
                           ALU_REG_out(28) => alu_out2_s_28_port, 
                           ALU_REG_out(27) => alu_out2_s_27_port, 
                           ALU_REG_out(26) => alu_out2_s_26_port, 
                           ALU_REG_out(25) => alu_out2_s_25_port, 
                           ALU_REG_out(24) => alu_out2_s_24_port, 
                           ALU_REG_out(23) => alu_out2_s_23_port, 
                           ALU_REG_out(22) => alu_out2_s_22_port, 
                           ALU_REG_out(21) => alu_out2_s_21_port, 
                           ALU_REG_out(20) => alu_out2_s_20_port, 
                           ALU_REG_out(19) => alu_out2_s_19_port, 
                           ALU_REG_out(18) => alu_out2_s_18_port, 
                           ALU_REG_out(17) => alu_out2_s_17_port, 
                           ALU_REG_out(16) => alu_out2_s_16_port, 
                           ALU_REG_out(15) => alu_out2_s_15_port, 
                           ALU_REG_out(14) => alu_out2_s_14_port, 
                           ALU_REG_out(13) => alu_out2_s_13_port, 
                           ALU_REG_out(12) => alu_out2_s_12_port, 
                           ALU_REG_out(11) => alu_out2_s_11_port, 
                           ALU_REG_out(10) => alu_out2_s_10_port, 
                           ALU_REG_out(9) => alu_out2_s_9_port, ALU_REG_out(8) 
                           => alu_out2_s_8_port, ALU_REG_out(7) => 
                           alu_out2_s_7_port, ALU_REG_out(6) => 
                           alu_out2_s_6_port, ALU_REG_out(5) => 
                           alu_out2_s_5_port, ALU_REG_out(4) => 
                           alu_out2_s_4_port, ALU_REG_out(3) => 
                           alu_out2_s_3_port, ALU_REG_out(2) => 
                           alu_out2_s_2_port, ALU_REG_out(1) => 
                           alu_out2_s_1_port, ALU_REG_out(0) => 
                           alu_out2_s_0_port, RT_REG_out(31) => 
                           rt_reg3_s_31_port, RT_REG_out(30) => 
                           rt_reg3_s_30_port, RT_REG_out(29) => 
                           rt_reg3_s_29_port, RT_REG_out(28) => 
                           rt_reg3_s_28_port, RT_REG_out(27) => 
                           rt_reg3_s_27_port, RT_REG_out(26) => 
                           rt_reg3_s_26_port, RT_REG_out(25) => 
                           rt_reg3_s_25_port, RT_REG_out(24) => 
                           rt_reg3_s_24_port, RT_REG_out(23) => 
                           rt_reg3_s_23_port, RT_REG_out(22) => 
                           rt_reg3_s_22_port, RT_REG_out(21) => 
                           rt_reg3_s_21_port, RT_REG_out(20) => 
                           rt_reg3_s_20_port, RT_REG_out(19) => 
                           rt_reg3_s_19_port, RT_REG_out(18) => 
                           rt_reg3_s_18_port, RT_REG_out(17) => 
                           rt_reg3_s_17_port, RT_REG_out(16) => 
                           rt_reg3_s_16_port, RT_REG_out(15) => 
                           rt_reg3_s_15_port, RT_REG_out(14) => 
                           rt_reg3_s_14_port, RT_REG_out(13) => 
                           rt_reg3_s_13_port, RT_REG_out(12) => 
                           rt_reg3_s_12_port, RT_REG_out(11) => 
                           rt_reg3_s_11_port, RT_REG_out(10) => 
                           rt_reg3_s_10_port, RT_REG_out(9) => rt_reg3_s_9_port
                           , RT_REG_out(8) => rt_reg3_s_8_port, RT_REG_out(7) 
                           => rt_reg3_s_7_port, RT_REG_out(6) => 
                           rt_reg3_s_6_port, RT_REG_out(5) => rt_reg3_s_5_port,
                           RT_REG_out(4) => rt_reg3_s_4_port, RT_REG_out(3) => 
                           rt_reg3_s_3_port, RT_REG_out(2) => rt_reg3_s_2_port,
                           RT_REG_out(1) => rt_reg3_s_1_port, RT_REG_out(0) => 
                           rt_reg3_s_0_port, NPC_REG_out(31) => 
                           npc_reg4_s_31_port, NPC_REG_out(30) => 
                           npc_reg4_s_30_port, NPC_REG_out(29) => 
                           npc_reg4_s_29_port, NPC_REG_out(28) => 
                           npc_reg4_s_28_port, NPC_REG_out(27) => 
                           npc_reg4_s_27_port, NPC_REG_out(26) => 
                           npc_reg4_s_26_port, NPC_REG_out(25) => 
                           npc_reg4_s_25_port, NPC_REG_out(24) => 
                           npc_reg4_s_24_port, NPC_REG_out(23) => 
                           npc_reg4_s_23_port, NPC_REG_out(22) => 
                           npc_reg4_s_22_port, NPC_REG_out(21) => 
                           npc_reg4_s_21_port, NPC_REG_out(20) => 
                           npc_reg4_s_20_port, NPC_REG_out(19) => 
                           npc_reg4_s_19_port, NPC_REG_out(18) => 
                           npc_reg4_s_18_port, NPC_REG_out(17) => 
                           npc_reg4_s_17_port, NPC_REG_out(16) => 
                           npc_reg4_s_16_port, NPC_REG_out(15) => 
                           npc_reg4_s_15_port, NPC_REG_out(14) => 
                           npc_reg4_s_14_port, NPC_REG_out(13) => 
                           npc_reg4_s_13_port, NPC_REG_out(12) => 
                           npc_reg4_s_12_port, NPC_REG_out(11) => 
                           npc_reg4_s_11_port, NPC_REG_out(10) => 
                           npc_reg4_s_10_port, NPC_REG_out(9) => 
                           npc_reg4_s_9_port, NPC_REG_out(8) => 
                           npc_reg4_s_8_port, NPC_REG_out(7) => 
                           npc_reg4_s_7_port, NPC_REG_out(6) => 
                           npc_reg4_s_6_port, NPC_REG_out(5) => 
                           npc_reg4_s_5_port, NPC_REG_out(4) => 
                           npc_reg4_s_4_port, NPC_REG_out(3) => 
                           npc_reg4_s_3_port, NPC_REG_out(2) => 
                           npc_reg4_s_2_port, NPC_REG_out(1) => 
                           npc_reg4_s_1_port, NPC_REG_out(0) => 
                           npc_reg4_s_0_port);
   WB_STAGE : WBU_N32 port map( ALU_OUT(31) => alu_out2_s_31_port, ALU_OUT(30) 
                           => alu_out2_s_30_port, ALU_OUT(29) => 
                           alu_out2_s_29_port, ALU_OUT(28) => 
                           alu_out2_s_28_port, ALU_OUT(27) => 
                           alu_out2_s_27_port, ALU_OUT(26) => 
                           alu_out2_s_26_port, ALU_OUT(25) => 
                           alu_out2_s_25_port, ALU_OUT(24) => 
                           alu_out2_s_24_port, ALU_OUT(23) => 
                           alu_out2_s_23_port, ALU_OUT(22) => 
                           alu_out2_s_22_port, ALU_OUT(21) => 
                           alu_out2_s_21_port, ALU_OUT(20) => 
                           alu_out2_s_20_port, ALU_OUT(19) => 
                           alu_out2_s_19_port, ALU_OUT(18) => 
                           alu_out2_s_18_port, ALU_OUT(17) => 
                           alu_out2_s_17_port, ALU_OUT(16) => 
                           alu_out2_s_16_port, ALU_OUT(15) => 
                           alu_out2_s_15_port, ALU_OUT(14) => 
                           alu_out2_s_14_port, ALU_OUT(13) => 
                           alu_out2_s_13_port, ALU_OUT(12) => 
                           alu_out2_s_12_port, ALU_OUT(11) => 
                           alu_out2_s_11_port, ALU_OUT(10) => 
                           alu_out2_s_10_port, ALU_OUT(9) => alu_out2_s_9_port,
                           ALU_OUT(8) => alu_out2_s_8_port, ALU_OUT(7) => 
                           alu_out2_s_7_port, ALU_OUT(6) => alu_out2_s_6_port, 
                           ALU_OUT(5) => alu_out2_s_5_port, ALU_OUT(4) => 
                           alu_out2_s_4_port, ALU_OUT(3) => alu_out2_s_3_port, 
                           ALU_OUT(2) => alu_out2_s_2_port, ALU_OUT(1) => 
                           alu_out2_s_1_port, ALU_OUT(0) => alu_out2_s_0_port, 
                           LOAD(31) => lmd_out_s_31_port, LOAD(30) => 
                           lmd_out_s_30_port, LOAD(29) => lmd_out_s_29_port, 
                           LOAD(28) => lmd_out_s_28_port, LOAD(27) => 
                           lmd_out_s_27_port, LOAD(26) => lmd_out_s_26_port, 
                           LOAD(25) => lmd_out_s_25_port, LOAD(24) => 
                           lmd_out_s_24_port, LOAD(23) => lmd_out_s_23_port, 
                           LOAD(22) => lmd_out_s_22_port, LOAD(21) => 
                           lmd_out_s_21_port, LOAD(20) => lmd_out_s_20_port, 
                           LOAD(19) => lmd_out_s_19_port, LOAD(18) => 
                           lmd_out_s_18_port, LOAD(17) => lmd_out_s_17_port, 
                           LOAD(16) => lmd_out_s_16_port, LOAD(15) => 
                           lmd_out_s_15_port, LOAD(14) => lmd_out_s_14_port, 
                           LOAD(13) => lmd_out_s_13_port, LOAD(12) => 
                           lmd_out_s_12_port, LOAD(11) => lmd_out_s_11_port, 
                           LOAD(10) => lmd_out_s_10_port, LOAD(9) => 
                           lmd_out_s_9_port, LOAD(8) => lmd_out_s_8_port, 
                           LOAD(7) => lmd_out_s_7_port, LOAD(6) => 
                           lmd_out_s_6_port, LOAD(5) => lmd_out_s_5_port, 
                           LOAD(4) => lmd_out_s_4_port, LOAD(3) => 
                           lmd_out_s_3_port, LOAD(2) => lmd_out_s_2_port, 
                           LOAD(1) => lmd_out_s_1_port, LOAD(0) => 
                           lmd_out_s_0_port, NPC_REG_in(31) => 
                           npc_reg4_s_31_port, NPC_REG_in(30) => 
                           npc_reg4_s_30_port, NPC_REG_in(29) => 
                           npc_reg4_s_29_port, NPC_REG_in(28) => 
                           npc_reg4_s_28_port, NPC_REG_in(27) => 
                           npc_reg4_s_27_port, NPC_REG_in(26) => 
                           npc_reg4_s_26_port, NPC_REG_in(25) => 
                           npc_reg4_s_25_port, NPC_REG_in(24) => 
                           npc_reg4_s_24_port, NPC_REG_in(23) => 
                           npc_reg4_s_23_port, NPC_REG_in(22) => 
                           npc_reg4_s_22_port, NPC_REG_in(21) => 
                           npc_reg4_s_21_port, NPC_REG_in(20) => 
                           npc_reg4_s_20_port, NPC_REG_in(19) => 
                           npc_reg4_s_19_port, NPC_REG_in(18) => 
                           npc_reg4_s_18_port, NPC_REG_in(17) => 
                           npc_reg4_s_17_port, NPC_REG_in(16) => 
                           npc_reg4_s_16_port, NPC_REG_in(15) => 
                           npc_reg4_s_15_port, NPC_REG_in(14) => 
                           npc_reg4_s_14_port, NPC_REG_in(13) => 
                           npc_reg4_s_13_port, NPC_REG_in(12) => 
                           npc_reg4_s_12_port, NPC_REG_in(11) => 
                           npc_reg4_s_11_port, NPC_REG_in(10) => 
                           npc_reg4_s_10_port, NPC_REG_in(9) => 
                           npc_reg4_s_9_port, NPC_REG_in(8) => 
                           npc_reg4_s_8_port, NPC_REG_in(7) => 
                           npc_reg4_s_7_port, NPC_REG_in(6) => 
                           npc_reg4_s_6_port, NPC_REG_in(5) => 
                           npc_reg4_s_5_port, NPC_REG_in(4) => 
                           npc_reg4_s_4_port, NPC_REG_in(3) => 
                           npc_reg4_s_3_port, NPC_REG_in(2) => 
                           npc_reg4_s_2_port, NPC_REG_in(1) => 
                           npc_reg4_s_1_port, NPC_REG_in(0) => 
                           npc_reg4_s_0_port, RT_REG_in(31) => 
                           rt_reg3_s_31_port, RT_REG_in(30) => 
                           rt_reg3_s_30_port, RT_REG_in(29) => 
                           rt_reg3_s_29_port, RT_REG_in(28) => 
                           rt_reg3_s_28_port, RT_REG_in(27) => 
                           rt_reg3_s_27_port, RT_REG_in(26) => 
                           rt_reg3_s_26_port, RT_REG_in(25) => 
                           rt_reg3_s_25_port, RT_REG_in(24) => 
                           rt_reg3_s_24_port, RT_REG_in(23) => 
                           rt_reg3_s_23_port, RT_REG_in(22) => 
                           rt_reg3_s_22_port, RT_REG_in(21) => 
                           rt_reg3_s_21_port, RT_REG_in(20) => 
                           rt_reg3_s_20_port, RT_REG_in(19) => 
                           rt_reg3_s_19_port, RT_REG_in(18) => 
                           rt_reg3_s_18_port, RT_REG_in(17) => 
                           rt_reg3_s_17_port, RT_REG_in(16) => 
                           rt_reg3_s_16_port, RT_REG_in(15) => 
                           rt_reg3_s_15_port, RT_REG_in(14) => 
                           rt_reg3_s_14_port, RT_REG_in(13) => 
                           rt_reg3_s_13_port, RT_REG_in(12) => 
                           rt_reg3_s_12_port, RT_REG_in(11) => 
                           rt_reg3_s_11_port, RT_REG_in(10) => 
                           rt_reg3_s_10_port, RT_REG_in(9) => rt_reg3_s_9_port,
                           RT_REG_in(8) => rt_reg3_s_8_port, RT_REG_in(7) => 
                           rt_reg3_s_7_port, RT_REG_in(6) => rt_reg3_s_6_port, 
                           RT_REG_in(5) => rt_reg3_s_5_port, RT_REG_in(4) => 
                           rt_reg3_s_4_port, RT_REG_in(3) => rt_reg3_s_3_port, 
                           RT_REG_in(2) => rt_reg3_s_2_port, RT_REG_in(1) => 
                           rt_reg3_s_1_port, RT_REG_in(0) => rt_reg3_s_0_port, 
                           IS_JAL => JAL_EN, ALUOUT_OR_LOAD => WB_MUX_SEL, 
                           RF_ADDR(31) => wb_addr_s_31_port, RF_ADDR(30) => 
                           wb_addr_s_30_port, RF_ADDR(29) => wb_addr_s_29_port,
                           RF_ADDR(28) => wb_addr_s_28_port, RF_ADDR(27) => 
                           wb_addr_s_27_port, RF_ADDR(26) => wb_addr_s_26_port,
                           RF_ADDR(25) => wb_addr_s_25_port, RF_ADDR(24) => 
                           wb_addr_s_24_port, RF_ADDR(23) => wb_addr_s_23_port,
                           RF_ADDR(22) => wb_addr_s_22_port, RF_ADDR(21) => 
                           wb_addr_s_21_port, RF_ADDR(20) => wb_addr_s_20_port,
                           RF_ADDR(19) => wb_addr_s_19_port, RF_ADDR(18) => 
                           wb_addr_s_18_port, RF_ADDR(17) => wb_addr_s_17_port,
                           RF_ADDR(16) => wb_addr_s_16_port, RF_ADDR(15) => 
                           wb_addr_s_15_port, RF_ADDR(14) => wb_addr_s_14_port,
                           RF_ADDR(13) => wb_addr_s_13_port, RF_ADDR(12) => 
                           wb_addr_s_12_port, RF_ADDR(11) => wb_addr_s_11_port,
                           RF_ADDR(10) => wb_addr_s_10_port, RF_ADDR(9) => 
                           wb_addr_s_9_port, RF_ADDR(8) => wb_addr_s_8_port, 
                           RF_ADDR(7) => wb_addr_s_7_port, RF_ADDR(6) => 
                           wb_addr_s_6_port, RF_ADDR(5) => wb_addr_s_5_port, 
                           RF_ADDR(4) => wb_addr_s_4_port, RF_ADDR(3) => 
                           wb_addr_s_3_port, RF_ADDR(2) => wb_addr_s_2_port, 
                           RF_ADDR(1) => wb_addr_s_1_port, RF_ADDR(0) => 
                           wb_addr_s_0_port, RF_DATA(31) => wb_data_s_31_port, 
                           RF_DATA(30) => wb_data_s_30_port, RF_DATA(29) => 
                           wb_data_s_29_port, RF_DATA(28) => wb_data_s_28_port,
                           RF_DATA(27) => wb_data_s_27_port, RF_DATA(26) => 
                           wb_data_s_26_port, RF_DATA(25) => wb_data_s_25_port,
                           RF_DATA(24) => wb_data_s_24_port, RF_DATA(23) => 
                           wb_data_s_23_port, RF_DATA(22) => wb_data_s_22_port,
                           RF_DATA(21) => wb_data_s_21_port, RF_DATA(20) => 
                           wb_data_s_20_port, RF_DATA(19) => wb_data_s_19_port,
                           RF_DATA(18) => wb_data_s_18_port, RF_DATA(17) => 
                           wb_data_s_17_port, RF_DATA(16) => wb_data_s_16_port,
                           RF_DATA(15) => wb_data_s_15_port, RF_DATA(14) => 
                           wb_data_s_14_port, RF_DATA(13) => wb_data_s_13_port,
                           RF_DATA(12) => wb_data_s_12_port, RF_DATA(11) => 
                           wb_data_s_11_port, RF_DATA(10) => wb_data_s_10_port,
                           RF_DATA(9) => wb_data_s_9_port, RF_DATA(8) => 
                           wb_data_s_8_port, RF_DATA(7) => wb_data_s_7_port, 
                           RF_DATA(6) => wb_data_s_6_port, RF_DATA(5) => 
                           wb_data_s_5_port, RF_DATA(4) => wb_data_s_4_port, 
                           RF_DATA(3) => wb_data_s_3_port, RF_DATA(2) => 
                           wb_data_s_2_port, RF_DATA(1) => wb_data_s_1_port, 
                           RF_DATA(0) => wb_data_s_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic;  DRAM_LMD, IRAM_IR : in std_logic_vector (31 
         downto 0);  DRAM_address, DRAM_data_in, IRAM_PC : out std_logic_vector
         (31 downto 0));

end DLX;

architecture SYN_dlx_rtl of DLX is

   component 
      dlx_cu_MICROCODE_MEM_SIZE33_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE19
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  branch_taken : in std_logic;  IR_EN, NPC_EN, RegA_EN, RegB_EN, 
            RegIMM_EN, RT_REG_EN, IS_R_TYPE, J_EN, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, BRANCH_EN, BEQZ_OR_BNEZ, SH2_EN : out std_logic;  
            ALU_OPCODE : out std_logic_vector (0 to 3);  DRAM_WE, LMD_EN, 
            WB_MUX_SEL, RF_WE, JAL_EN, PC_EN : out std_logic);
   end component;
   
   component DATAPATH_N32
      port( CLK, RST : in std_logic;  ALU_FUNC : in std_logic_vector (0 to 3); 
            from_IRAM, from_DRAM : in std_logic_vector (31 downto 0);  IR_EN, 
            NPC_EN, RegA_EN, RegB_EN, RegIMM_EN, RT_REG_EN, IS_R_TYPE, J_EN, 
            MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, BRANCH_EN, BEQZ_OR_BNEZ, SH2_EN,
            LMD_EN, WB_MUX_SEL, RF_WE, JAL_EN, PC_EN : in std_logic;  
            branch_taken : out std_logic;  addr_to_DRAM, data_to_DRAM, to_IRAM,
            IR : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, ALU_OPCODE_i_0_port, ALU_OPCODE_i_1_port, 
      ALU_OPCODE_i_2_port, ALU_OPCODE_i_3_port, IR_EN_i, NPC_EN_i, RegA_EN_i, 
      RegB_EN_i, RegIMM_EN_i, RT_REG_EN_i, IS_R_TYPE_i, J_EN_i, MUXA_SEL_i, 
      MUXB_SEL_i, ALU_OUTREG_EN_i, BEQZ_OR_BNEZ_i, SH2_EN_i, LMD_EN_i, 
      WB_MUX_SEL_i, RF_WE_i, JAL_EN_i, PC_EN_i, branch_taken_i, n_1673, n_1674,
      n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, 
      n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, 
      n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, 
      n_1702, n_1703, n_1704, n_1705, n_1706, n_1707 : std_logic;

begin
   
   X_Logic0_port <= '0';
   PC_EN_i <= '1';
   DATAPATH_I : DATAPATH_N32 port map( CLK => Clk, RST => Rst, ALU_FUNC(0) => 
                           ALU_OPCODE_i_0_port, ALU_FUNC(1) => 
                           ALU_OPCODE_i_1_port, ALU_FUNC(2) => 
                           ALU_OPCODE_i_2_port, ALU_FUNC(3) => 
                           ALU_OPCODE_i_3_port, from_IRAM(31) => IRAM_IR(31), 
                           from_IRAM(30) => IRAM_IR(30), from_IRAM(29) => 
                           IRAM_IR(29), from_IRAM(28) => IRAM_IR(28), 
                           from_IRAM(27) => IRAM_IR(27), from_IRAM(26) => 
                           IRAM_IR(26), from_IRAM(25) => IRAM_IR(25), 
                           from_IRAM(24) => IRAM_IR(24), from_IRAM(23) => 
                           IRAM_IR(23), from_IRAM(22) => IRAM_IR(22), 
                           from_IRAM(21) => IRAM_IR(21), from_IRAM(20) => 
                           IRAM_IR(20), from_IRAM(19) => IRAM_IR(19), 
                           from_IRAM(18) => IRAM_IR(18), from_IRAM(17) => 
                           IRAM_IR(17), from_IRAM(16) => IRAM_IR(16), 
                           from_IRAM(15) => IRAM_IR(15), from_IRAM(14) => 
                           IRAM_IR(14), from_IRAM(13) => IRAM_IR(13), 
                           from_IRAM(12) => IRAM_IR(12), from_IRAM(11) => 
                           IRAM_IR(11), from_IRAM(10) => IRAM_IR(10), 
                           from_IRAM(9) => IRAM_IR(9), from_IRAM(8) => 
                           IRAM_IR(8), from_IRAM(7) => IRAM_IR(7), from_IRAM(6)
                           => IRAM_IR(6), from_IRAM(5) => IRAM_IR(5), 
                           from_IRAM(4) => IRAM_IR(4), from_IRAM(3) => 
                           IRAM_IR(3), from_IRAM(2) => IRAM_IR(2), from_IRAM(1)
                           => IRAM_IR(1), from_IRAM(0) => IRAM_IR(0), 
                           from_DRAM(31) => DRAM_LMD(31), from_DRAM(30) => 
                           DRAM_LMD(30), from_DRAM(29) => DRAM_LMD(29), 
                           from_DRAM(28) => DRAM_LMD(28), from_DRAM(27) => 
                           DRAM_LMD(27), from_DRAM(26) => DRAM_LMD(26), 
                           from_DRAM(25) => DRAM_LMD(25), from_DRAM(24) => 
                           DRAM_LMD(24), from_DRAM(23) => DRAM_LMD(23), 
                           from_DRAM(22) => DRAM_LMD(22), from_DRAM(21) => 
                           DRAM_LMD(21), from_DRAM(20) => DRAM_LMD(20), 
                           from_DRAM(19) => DRAM_LMD(19), from_DRAM(18) => 
                           DRAM_LMD(18), from_DRAM(17) => DRAM_LMD(17), 
                           from_DRAM(16) => DRAM_LMD(16), from_DRAM(15) => 
                           DRAM_LMD(15), from_DRAM(14) => DRAM_LMD(14), 
                           from_DRAM(13) => DRAM_LMD(13), from_DRAM(12) => 
                           DRAM_LMD(12), from_DRAM(11) => DRAM_LMD(11), 
                           from_DRAM(10) => DRAM_LMD(10), from_DRAM(9) => 
                           DRAM_LMD(9), from_DRAM(8) => DRAM_LMD(8), 
                           from_DRAM(7) => DRAM_LMD(7), from_DRAM(6) => 
                           DRAM_LMD(6), from_DRAM(5) => DRAM_LMD(5), 
                           from_DRAM(4) => DRAM_LMD(4), from_DRAM(3) => 
                           DRAM_LMD(3), from_DRAM(2) => DRAM_LMD(2), 
                           from_DRAM(1) => DRAM_LMD(1), from_DRAM(0) => 
                           DRAM_LMD(0), IR_EN => IR_EN_i, NPC_EN => NPC_EN_i, 
                           RegA_EN => RegA_EN_i, RegB_EN => RegB_EN_i, 
                           RegIMM_EN => RegIMM_EN_i, RT_REG_EN => RT_REG_EN_i, 
                           IS_R_TYPE => IS_R_TYPE_i, J_EN => J_EN_i, MUXA_SEL 
                           => MUXA_SEL_i, MUXB_SEL => MUXB_SEL_i, ALU_OUTREG_EN
                           => ALU_OUTREG_EN_i, BRANCH_EN => X_Logic0_port, 
                           BEQZ_OR_BNEZ => BEQZ_OR_BNEZ_i, SH2_EN => SH2_EN_i, 
                           LMD_EN => LMD_EN_i, WB_MUX_SEL => WB_MUX_SEL_i, 
                           RF_WE => RF_WE_i, JAL_EN => JAL_EN_i, PC_EN => 
                           PC_EN_i, branch_taken => branch_taken_i, 
                           addr_to_DRAM(31) => DRAM_address(31), 
                           addr_to_DRAM(30) => DRAM_address(30), 
                           addr_to_DRAM(29) => DRAM_address(29), 
                           addr_to_DRAM(28) => DRAM_address(28), 
                           addr_to_DRAM(27) => DRAM_address(27), 
                           addr_to_DRAM(26) => DRAM_address(26), 
                           addr_to_DRAM(25) => DRAM_address(25), 
                           addr_to_DRAM(24) => DRAM_address(24), 
                           addr_to_DRAM(23) => DRAM_address(23), 
                           addr_to_DRAM(22) => DRAM_address(22), 
                           addr_to_DRAM(21) => DRAM_address(21), 
                           addr_to_DRAM(20) => DRAM_address(20), 
                           addr_to_DRAM(19) => DRAM_address(19), 
                           addr_to_DRAM(18) => DRAM_address(18), 
                           addr_to_DRAM(17) => DRAM_address(17), 
                           addr_to_DRAM(16) => DRAM_address(16), 
                           addr_to_DRAM(15) => DRAM_address(15), 
                           addr_to_DRAM(14) => DRAM_address(14), 
                           addr_to_DRAM(13) => DRAM_address(13), 
                           addr_to_DRAM(12) => DRAM_address(12), 
                           addr_to_DRAM(11) => DRAM_address(11), 
                           addr_to_DRAM(10) => DRAM_address(10), 
                           addr_to_DRAM(9) => DRAM_address(9), addr_to_DRAM(8) 
                           => DRAM_address(8), addr_to_DRAM(7) => 
                           DRAM_address(7), addr_to_DRAM(6) => DRAM_address(6),
                           addr_to_DRAM(5) => DRAM_address(5), addr_to_DRAM(4) 
                           => DRAM_address(4), addr_to_DRAM(3) => 
                           DRAM_address(3), addr_to_DRAM(2) => DRAM_address(2),
                           addr_to_DRAM(1) => DRAM_address(1), addr_to_DRAM(0) 
                           => DRAM_address(0), data_to_DRAM(31) => 
                           DRAM_data_in(31), data_to_DRAM(30) => 
                           DRAM_data_in(30), data_to_DRAM(29) => 
                           DRAM_data_in(29), data_to_DRAM(28) => 
                           DRAM_data_in(28), data_to_DRAM(27) => 
                           DRAM_data_in(27), data_to_DRAM(26) => 
                           DRAM_data_in(26), data_to_DRAM(25) => 
                           DRAM_data_in(25), data_to_DRAM(24) => 
                           DRAM_data_in(24), data_to_DRAM(23) => 
                           DRAM_data_in(23), data_to_DRAM(22) => 
                           DRAM_data_in(22), data_to_DRAM(21) => 
                           DRAM_data_in(21), data_to_DRAM(20) => 
                           DRAM_data_in(20), data_to_DRAM(19) => 
                           DRAM_data_in(19), data_to_DRAM(18) => 
                           DRAM_data_in(18), data_to_DRAM(17) => 
                           DRAM_data_in(17), data_to_DRAM(16) => 
                           DRAM_data_in(16), data_to_DRAM(15) => 
                           DRAM_data_in(15), data_to_DRAM(14) => 
                           DRAM_data_in(14), data_to_DRAM(13) => 
                           DRAM_data_in(13), data_to_DRAM(12) => 
                           DRAM_data_in(12), data_to_DRAM(11) => 
                           DRAM_data_in(11), data_to_DRAM(10) => 
                           DRAM_data_in(10), data_to_DRAM(9) => DRAM_data_in(9)
                           , data_to_DRAM(8) => DRAM_data_in(8), 
                           data_to_DRAM(7) => DRAM_data_in(7), data_to_DRAM(6) 
                           => DRAM_data_in(6), data_to_DRAM(5) => 
                           DRAM_data_in(5), data_to_DRAM(4) => DRAM_data_in(4),
                           data_to_DRAM(3) => DRAM_data_in(3), data_to_DRAM(2) 
                           => DRAM_data_in(2), data_to_DRAM(1) => 
                           DRAM_data_in(1), data_to_DRAM(0) => DRAM_data_in(0),
                           to_IRAM(31) => IRAM_PC(31), to_IRAM(30) => 
                           IRAM_PC(30), to_IRAM(29) => IRAM_PC(29), to_IRAM(28)
                           => IRAM_PC(28), to_IRAM(27) => IRAM_PC(27), 
                           to_IRAM(26) => IRAM_PC(26), to_IRAM(25) => 
                           IRAM_PC(25), to_IRAM(24) => IRAM_PC(24), to_IRAM(23)
                           => IRAM_PC(23), to_IRAM(22) => IRAM_PC(22), 
                           to_IRAM(21) => IRAM_PC(21), to_IRAM(20) => 
                           IRAM_PC(20), to_IRAM(19) => IRAM_PC(19), to_IRAM(18)
                           => IRAM_PC(18), to_IRAM(17) => IRAM_PC(17), 
                           to_IRAM(16) => IRAM_PC(16), to_IRAM(15) => 
                           IRAM_PC(15), to_IRAM(14) => IRAM_PC(14), to_IRAM(13)
                           => IRAM_PC(13), to_IRAM(12) => IRAM_PC(12), 
                           to_IRAM(11) => IRAM_PC(11), to_IRAM(10) => 
                           IRAM_PC(10), to_IRAM(9) => IRAM_PC(9), to_IRAM(8) =>
                           IRAM_PC(8), to_IRAM(7) => IRAM_PC(7), to_IRAM(6) => 
                           IRAM_PC(6), to_IRAM(5) => IRAM_PC(5), to_IRAM(4) => 
                           IRAM_PC(4), to_IRAM(3) => IRAM_PC(3), to_IRAM(2) => 
                           IRAM_PC(2), to_IRAM(1) => IRAM_PC(1), to_IRAM(0) => 
                           IRAM_PC(0), IR(31) => n_1673, IR(30) => n_1674, 
                           IR(29) => n_1675, IR(28) => n_1676, IR(27) => n_1677
                           , IR(26) => n_1678, IR(25) => n_1679, IR(24) => 
                           n_1680, IR(23) => n_1681, IR(22) => n_1682, IR(21) 
                           => n_1683, IR(20) => n_1684, IR(19) => n_1685, 
                           IR(18) => n_1686, IR(17) => n_1687, IR(16) => n_1688
                           , IR(15) => n_1689, IR(14) => n_1690, IR(13) => 
                           n_1691, IR(12) => n_1692, IR(11) => n_1693, IR(10) 
                           => n_1694, IR(9) => n_1695, IR(8) => n_1696, IR(7) 
                           => n_1697, IR(6) => n_1698, IR(5) => n_1699, IR(4) 
                           => n_1700, IR(3) => n_1701, IR(2) => n_1702, IR(1) 
                           => n_1703, IR(0) => n_1704);
   CU_I : 
                           dlx_cu_MICROCODE_MEM_SIZE33_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE19 
                           port map( Clk => Clk, Rst => Rst, IR_IN(31) => 
                           IRAM_IR(31), IR_IN(30) => IRAM_IR(30), IR_IN(29) => 
                           IRAM_IR(29), IR_IN(28) => IRAM_IR(28), IR_IN(27) => 
                           IRAM_IR(27), IR_IN(26) => IRAM_IR(26), IR_IN(25) => 
                           IRAM_IR(25), IR_IN(24) => IRAM_IR(24), IR_IN(23) => 
                           IRAM_IR(23), IR_IN(22) => IRAM_IR(22), IR_IN(21) => 
                           IRAM_IR(21), IR_IN(20) => IRAM_IR(20), IR_IN(19) => 
                           IRAM_IR(19), IR_IN(18) => IRAM_IR(18), IR_IN(17) => 
                           IRAM_IR(17), IR_IN(16) => IRAM_IR(16), IR_IN(15) => 
                           IRAM_IR(15), IR_IN(14) => IRAM_IR(14), IR_IN(13) => 
                           IRAM_IR(13), IR_IN(12) => IRAM_IR(12), IR_IN(11) => 
                           IRAM_IR(11), IR_IN(10) => IRAM_IR(10), IR_IN(9) => 
                           IRAM_IR(9), IR_IN(8) => IRAM_IR(8), IR_IN(7) => 
                           IRAM_IR(7), IR_IN(6) => IRAM_IR(6), IR_IN(5) => 
                           IRAM_IR(5), IR_IN(4) => IRAM_IR(4), IR_IN(3) => 
                           IRAM_IR(3), IR_IN(2) => IRAM_IR(2), IR_IN(1) => 
                           IRAM_IR(1), IR_IN(0) => IRAM_IR(0), branch_taken => 
                           branch_taken_i, IR_EN => IR_EN_i, NPC_EN => NPC_EN_i
                           , RegA_EN => RegA_EN_i, RegB_EN => RegB_EN_i, 
                           RegIMM_EN => RegIMM_EN_i, RT_REG_EN => RT_REG_EN_i, 
                           IS_R_TYPE => IS_R_TYPE_i, J_EN => J_EN_i, MUXA_SEL 
                           => MUXA_SEL_i, MUXB_SEL => MUXB_SEL_i, ALU_OUTREG_EN
                           => ALU_OUTREG_EN_i, BRANCH_EN => n_1705, 
                           BEQZ_OR_BNEZ => BEQZ_OR_BNEZ_i, SH2_EN => SH2_EN_i, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_0_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_1_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_3_port, DRAM_WE => n_1706, LMD_EN => 
                           LMD_EN_i, WB_MUX_SEL => WB_MUX_SEL_i, RF_WE => 
                           RF_WE_i, JAL_EN => JAL_EN_i, PC_EN => n_1707);

end SYN_dlx_rtl;
